-- x49_shares
-- Input_shares: X00, X0_1, X02, X03; X10, X11, X12, X13; X20, X21, X22, X23; X30, X31, X32, X33; X40, X41, X42, X43; X50, X51, X52, X53; X60, X61, X62, X63; X70, X71, X72, X73.
-- Output_shares: F00, F01, F02, F03; F10, F11, F12, F13; F20, F21, F22, F23; F30, F31, F32, F33; F40, F41, F42, F43; F50, F51, F52, F53; F60, F61, F62, F63; F70, F71, F72, F73.
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity x49_shares is
    port (
    X00, X0_1, X02, X03, X10, X11, X12, X13, X20, X21, X22, X23, X30, X31, X32, X33, X40, X41, X42, X43, X50, X51, X52, X53, X60, X61, X62, X63, X70, X71, X72, X73 : in std_logic;
    F00, F01, F02, F03, F10, F11, F12, F13, F20, F21, F22, F23, F30, F31, F32, F33, F40, F41, F42, F43, F50, F51, F52, F53, F60, F61, F62, F63, F70, F71, F72, F73 : out std_logic);
end x49_shares;
architecture Behavioral of x49_shares is
begin
    F00  <= ((X00) xor (X10) xor (X00 and X10) xor (X00 and X11) xor (X02 and X10) xor (X00 and X12) xor (X10 and X20) xor (X10 and X21) xor (X12 and X20) xor (X10 and X22) xor (X00 and X10 and X20) xor (X00 and X10 and X22) xor (X00 and X11 and X21) xor (X00 and X11 and X22) xor (X00 and X12 and X21) xor (X0_1 and X10 and X20) xor (X0_1 and X10 and X22) xor (X0_1 and X11 and X20) xor (X0_1 and X12 and X20) xor (X0_1 and X12 and X21) xor (X02 and X10 and X20) xor (X02 and X10 and X21) xor (X02 and X11 and X20) xor (X02 and X11 and X21) xor (X02 and X12 and X20) xor (X02 and X12 and X22) xor (X30) xor (X10 and X30) xor (X10 and X31) xor (X12 and X30) xor (X10 and X32) xor (X00 and X10 and X30) xor (X00 and X10 and X32) xor (X00 and X11 and X31) xor (X00 and X11 and X32) xor (X00 and X12 and X31) xor (X0_1 and X10 and X30) xor (X0_1 and X10 and X32) xor (X0_1 and X11 and X30) xor (X0_1 and X12 and X30) xor (X0_1 and X12 and X31) xor (X02 and X10 and X30) xor (X02 and X10 and X31) xor (X02 and X11 and X30) xor (X02 and X11 and X31) xor (X02 and X12 and X30) xor (X02 and X12 and X32) xor (X20 and X30) xor (X20 and X31) xor (X22 and X30) xor (X20 and X32) xor (X10 and X40) xor (X10 and X41) xor (X12 and X40) xor (X10 and X42) xor (X00 and X10 and X40) xor (X00 and X10 and X42) xor (X00 and X11 and X41) xor (X00 and X11 and X42) xor (X00 and X12 and X41) xor (X0_1 and X10 and X40) xor (X0_1 and X10 and X42) xor (X0_1 and X11 and X40) xor (X0_1 and X12 and X40) xor (X0_1 and X12 and X41) xor (X02 and X10 and X40) xor (X02 and X10 and X41) xor (X02 and X11 and X40) xor (X02 and X11 and X41) xor (X02 and X12 and X40) xor (X02 and X12 and X42) xor (X30 and X40) xor (X30 and X41) xor (X32 and X40) xor (X30 and X42) xor (X20 and X30 and X40) xor (X20 and X30 and X42) xor (X20 and X31 and X41) xor (X20 and X31 and X42) xor (X20 and X32 and X41) xor (X21 and X30 and X40) xor (X21 and X30 and X42) xor (X21 and X31 and X40) xor (X21 and X32 and X40) xor (X21 and X32 and X41) xor (X22 and X30 and X40) xor (X22 and X30 and X41) xor (X22 and X31 and X40) xor (X22 and X31 and X41) xor (X22 and X32 and X40) xor (X22 and X32 and X42) xor (X50) xor (X00 and X50) xor (X00 and X51) xor (X02 and X50) xor (X00 and X52) xor (X20 and X50) xor (X20 and X51) xor (X22 and X50) xor (X20 and X52) xor (X30 and X50) xor (X30 and X51) xor (X32 and X50) xor (X30 and X52) xor (X00 and X30 and X50) xor (X00 and X30 and X52) xor (X00 and X31 and X51) xor (X00 and X31 and X52) xor (X00 and X32 and X51) xor (X0_1 and X30 and X50) xor (X0_1 and X30 and X52) xor (X0_1 and X31 and X50) xor (X0_1 and X32 and X50) xor (X0_1 and X32 and X51) xor (X02 and X30 and X50) xor (X02 and X30 and X51) xor (X02 and X31 and X50) xor (X02 and X31 and X51) xor (X02 and X32 and X50) xor (X02 and X32 and X52) xor (X20 and X30 and X50) xor (X20 and X30 and X52) xor (X20 and X31 and X51) xor (X20 and X31 and X52) xor (X20 and X32 and X51) xor (X21 and X30 and X50) xor (X21 and X30 and X52) xor (X21 and X31 and X50) xor (X21 and X32 and X50) xor (X21 and X32 and X51) xor (X22 and X30 and X50) xor (X22 and X30 and X51) xor (X22 and X31 and X50) xor (X22 and X31 and X51) xor (X22 and X32 and X50) xor (X22 and X32 and X52) xor (X00 and X40 and X50) xor (X00 and X40 and X52) xor (X00 and X41 and X51) xor (X00 and X41 and X52) xor (X00 and X42 and X51) xor (X0_1 and X40 and X50) xor (X0_1 and X40 and X52) xor (X0_1 and X41 and X50) xor (X0_1 and X42 and X50) xor (X0_1 and X42 and X51) xor (X02 and X40 and X50) xor (X02 and X40 and X51) xor (X02 and X41 and X50) xor (X02 and X41 and X51) xor (X02 and X42 and X50) xor (X02 and X42 and X52) xor (X10 and X40 and X50) xor (X10 and X40 and X52) xor (X10 and X41 and X51) xor (X10 and X41 and X52) xor (X10 and X42 and X51) xor (X11 and X40 and X50) xor (X11 and X40 and X52) xor (X11 and X41 and X50) xor (X11 and X42 and X50) xor (X11 and X42 and X51) xor (X12 and X40 and X50) xor (X12 and X40 and X51) xor (X12 and X41 and X50) xor (X12 and X41 and X51) xor (X12 and X42 and X50) xor (X12 and X42 and X52) xor (X20 and X40 and X50) xor (X20 and X40 and X52) xor (X20 and X41 and X51) xor (X20 and X41 and X52) xor (X20 and X42 and X51) xor (X21 and X40 and X50) xor (X21 and X40 and X52) xor (X21 and X41 and X50) xor (X21 and X42 and X50) xor (X21 and X42 and X51) xor (X22 and X40 and X50) xor (X22 and X40 and X51) xor (X22 and X41 and X50) xor (X22 and X41 and X51) xor (X22 and X42 and X50) xor (X22 and X42 and X52) xor (X00 and X10 and X60) xor (X00 and X10 and X62) xor (X00 and X11 and X61) xor (X00 and X11 and X62) xor (X00 and X12 and X61) xor (X0_1 and X10 and X60) xor (X0_1 and X10 and X62) xor (X0_1 and X11 and X60) xor (X0_1 and X12 and X60) xor (X0_1 and X12 and X61) xor (X02 and X10 and X60) xor (X02 and X10 and X61) xor (X02 and X11 and X60) xor (X02 and X11 and X61) xor (X02 and X12 and X60) xor (X02 and X12 and X62) xor (X20 and X60) xor (X20 and X61) xor (X22 and X60) xor (X20 and X62) xor (X00 and X20 and X60) xor (X00 and X20 and X62) xor (X00 and X21 and X61) xor (X00 and X21 and X62) xor (X00 and X22 and X61) xor (X0_1 and X20 and X60) xor (X0_1 and X20 and X62) xor (X0_1 and X21 and X60) xor (X0_1 and X22 and X60) xor (X0_1 and X22 and X61) xor (X02 and X20 and X60) xor (X02 and X20 and X61) xor (X02 and X21 and X60) xor (X02 and X21 and X61) xor (X02 and X22 and X60) xor (X02 and X22 and X62) xor (X30 and X60) xor (X30 and X61) xor (X32 and X60) xor (X30 and X62) xor (X00 and X30 and X60) xor (X00 and X30 and X62) xor (X00 and X31 and X61) xor (X00 and X31 and X62) xor (X00 and X32 and X61) xor (X0_1 and X30 and X60) xor (X0_1 and X30 and X62) xor (X0_1 and X31 and X60) xor (X0_1 and X32 and X60) xor (X0_1 and X32 and X61) xor (X02 and X30 and X60) xor (X02 and X30 and X61) xor (X02 and X31 and X60) xor (X02 and X31 and X61) xor (X02 and X32 and X60) xor (X02 and X32 and X62) xor (X10 and X30 and X60) xor (X10 and X30 and X62) xor (X10 and X31 and X61) xor (X10 and X31 and X62) xor (X10 and X32 and X61) xor (X11 and X30 and X60) xor (X11 and X30 and X62) xor (X11 and X31 and X60) xor (X11 and X32 and X60) xor (X11 and X32 and X61) xor (X12 and X30 and X60) xor (X12 and X30 and X61) xor (X12 and X31 and X60) xor (X12 and X31 and X61) xor (X12 and X32 and X60) xor (X12 and X32 and X62) xor (X40 and X60) xor (X40 and X61) xor (X42 and X60) xor (X40 and X62) xor (X50 and X60) xor (X50 and X61) xor (X52 and X60) xor (X50 and X62) xor (X20 and X50 and X60) xor (X20 and X50 and X62) xor (X20 and X51 and X61) xor (X20 and X51 and X62) xor (X20 and X52 and X61) xor (X21 and X50 and X60) xor (X21 and X50 and X62) xor (X21 and X51 and X60) xor (X21 and X52 and X60) xor (X21 and X52 and X61) xor (X22 and X50 and X60) xor (X22 and X50 and X61) xor (X22 and X51 and X60) xor (X22 and X51 and X61) xor (X22 and X52 and X60) xor (X22 and X52 and X62) xor (X70) xor (X00 and X70) xor (X00 and X71) xor (X02 and X70) xor (X00 and X72) xor (X00 and X10 and X70) xor (X00 and X10 and X72) xor (X00 and X11 and X71) xor (X00 and X11 and X72) xor (X00 and X12 and X71) xor (X0_1 and X10 and X70) xor (X0_1 and X10 and X72) xor (X0_1 and X11 and X70) xor (X0_1 and X12 and X70) xor (X0_1 and X12 and X71) xor (X02 and X10 and X70) xor (X02 and X10 and X71) xor (X02 and X11 and X70) xor (X02 and X11 and X71) xor (X02 and X12 and X70) xor (X02 and X12 and X72) xor (X20 and X70) xor (X20 and X71) xor (X22 and X70) xor (X20 and X72) xor (X00 and X30 and X70) xor (X00 and X30 and X72) xor (X00 and X31 and X71) xor (X00 and X31 and X72) xor (X00 and X32 and X71) xor (X0_1 and X30 and X70) xor (X0_1 and X30 and X72) xor (X0_1 and X31 and X70) xor (X0_1 and X32 and X70) xor (X0_1 and X32 and X71) xor (X02 and X30 and X70) xor (X02 and X30 and X71) xor (X02 and X31 and X70) xor (X02 and X31 and X71) xor (X02 and X32 and X70) xor (X02 and X32 and X72) xor (X20 and X30 and X70) xor (X20 and X30 and X72) xor (X20 and X31 and X71) xor (X20 and X31 and X72) xor (X20 and X32 and X71) xor (X21 and X30 and X70) xor (X21 and X30 and X72) xor (X21 and X31 and X70) xor (X21 and X32 and X70) xor (X21 and X32 and X71) xor (X22 and X30 and X70) xor (X22 and X30 and X71) xor (X22 and X31 and X70) xor (X22 and X31 and X71) xor (X22 and X32 and X70) xor (X22 and X32 and X72) xor (X10 and X40 and X70) xor (X10 and X40 and X72) xor (X10 and X41 and X71) xor (X10 and X41 and X72) xor (X10 and X42 and X71) xor (X11 and X40 and X70) xor (X11 and X40 and X72) xor (X11 and X41 and X70) xor (X11 and X42 and X70) xor (X11 and X42 and X71) xor (X12 and X40 and X70) xor (X12 and X40 and X71) xor (X12 and X41 and X70) xor (X12 and X41 and X71) xor (X12 and X42 and X70) xor (X12 and X42 and X72) xor (X30 and X40 and X70) xor (X30 and X40 and X72) xor (X30 and X41 and X71) xor (X30 and X41 and X72) xor (X30 and X42 and X71) xor (X31 and X40 and X70) xor (X31 and X40 and X72) xor (X31 and X41 and X70) xor (X31 and X42 and X70) xor (X31 and X42 and X71) xor (X32 and X40 and X70) xor (X32 and X40 and X71) xor (X32 and X41 and X70) xor (X32 and X41 and X71) xor (X32 and X42 and X70) xor (X32 and X42 and X72) xor (X00 and X50 and X70) xor (X00 and X50 and X72) xor (X00 and X51 and X71) xor (X00 and X51 and X72) xor (X00 and X52 and X71) xor (X0_1 and X50 and X70) xor (X0_1 and X50 and X72) xor (X0_1 and X51 and X70) xor (X0_1 and X52 and X70) xor (X0_1 and X52 and X71) xor (X02 and X50 and X70) xor (X02 and X50 and X71) xor (X02 and X51 and X70) xor (X02 and X51 and X71) xor (X02 and X52 and X70) xor (X02 and X52 and X72) xor (X20 and X50 and X70) xor (X20 and X50 and X72) xor (X20 and X51 and X71) xor (X20 and X51 and X72) xor (X20 and X52 and X71) xor (X21 and X50 and X70) xor (X21 and X50 and X72) xor (X21 and X51 and X70) xor (X21 and X52 and X70) xor (X21 and X52 and X71) xor (X22 and X50 and X70) xor (X22 and X50 and X71) xor (X22 and X51 and X70) xor (X22 and X51 and X71) xor (X22 and X52 and X70) xor (X22 and X52 and X72) xor (X00 and X60 and X70) xor (X00 and X60 and X72) xor (X00 and X61 and X71) xor (X00 and X61 and X72) xor (X00 and X62 and X71) xor (X0_1 and X60 and X70) xor (X0_1 and X60 and X72) xor (X0_1 and X61 and X70) xor (X0_1 and X62 and X70) xor (X0_1 and X62 and X71) xor (X02 and X60 and X70) xor (X02 and X60 and X71) xor (X02 and X61 and X70) xor (X02 and X61 and X71) xor (X02 and X62 and X70) xor (X02 and X62 and X72) xor (X10 and X60 and X70) xor (X10 and X60 and X72) xor (X10 and X61 and X71) xor (X10 and X61 and X72) xor (X10 and X62 and X71) xor (X11 and X60 and X70) xor (X11 and X60 and X72) xor (X11 and X61 and X70) xor (X11 and X62 and X70) xor (X11 and X62 and X71) xor (X12 and X60 and X70) xor (X12 and X60 and X71) xor (X12 and X61 and X70) xor (X12 and X61 and X71) xor (X12 and X62 and X70) xor (X12 and X62 and X72) xor (X20 and X60 and X70) xor (X20 and X60 and X72) xor (X20 and X61 and X71) xor (X20 and X61 and X72) xor (X20 and X62 and X71) xor (X21 and X60 and X70) xor (X21 and X60 and X72) xor (X21 and X61 and X70) xor (X21 and X62 and X70) xor (X21 and X62 and X71) xor (X22 and X60 and X70) xor (X22 and X60 and X71) xor (X22 and X61 and X70) xor (X22 and X61 and X71) xor (X22 and X62 and X70) xor (X22 and X62 and X72) xor (X40 and X60 and X70) xor (X40 and X60 and X72) xor (X40 and X61 and X71) xor (X40 and X61 and X72) xor (X40 and X62 and X71) xor (X41 and X60 and X70) xor (X41 and X60 and X72) xor (X41 and X61 and X70) xor (X41 and X62 and X70) xor (X41 and X62 and X71) xor (X42 and X60 and X70) xor (X42 and X60 and X71) xor (X42 and X61 and X70) xor (X42 and X61 and X71) xor (X42 and X62 and X70) xor (X42 and X62 and X72));
    F01  <= ((X0_1) xor (X11) xor (X0_1 and X11) xor (X0_1 and X12) xor (X02 and X11) xor (X0_1 and X13) xor (X11 and X21) xor (X11 and X22) xor (X12 and X21) xor (X11 and X23) xor (X0_1 and X11 and X21) xor (X0_1 and X11 and X22) xor (X0_1 and X12 and X22) xor (X0_1 and X12 and X23) xor (X0_1 and X13 and X22) xor (X02 and X11 and X22) xor (X02 and X11 and X23) xor (X02 and X12 and X21) xor (X02 and X12 and X23) xor (X02 and X13 and X21) xor (X02 and X13 and X22) xor (X03 and X11 and X22) xor (X03 and X12 and X21) xor (X03 and X12 and X23) xor (X03 and X13 and X21) xor (X03 and X13 and X23) xor (X31) xor (X11 and X31) xor (X11 and X32) xor (X12 and X31) xor (X11 and X33) xor (X0_1 and X11 and X31) xor (X0_1 and X11 and X32) xor (X0_1 and X12 and X32) xor (X0_1 and X12 and X33) xor (X0_1 and X13 and X32) xor (X02 and X11 and X32) xor (X02 and X11 and X33) xor (X02 and X12 and X31) xor (X02 and X12 and X33) xor (X02 and X13 and X31) xor (X02 and X13 and X32) xor (X03 and X11 and X32) xor (X03 and X12 and X31) xor (X03 and X12 and X33) xor (X03 and X13 and X31) xor (X03 and X13 and X33) xor (X21 and X31) xor (X21 and X32) xor (X22 and X31) xor (X21 and X33) xor (X11 and X41) xor (X11 and X42) xor (X12 and X41) xor (X11 and X43) xor (X0_1 and X11 and X41) xor (X0_1 and X11 and X42) xor (X0_1 and X12 and X42) xor (X0_1 and X12 and X43) xor (X0_1 and X13 and X42) xor (X02 and X11 and X42) xor (X02 and X11 and X43) xor (X02 and X12 and X41) xor (X02 and X12 and X43) xor (X02 and X13 and X41) xor (X02 and X13 and X42) xor (X03 and X11 and X42) xor (X03 and X12 and X41) xor (X03 and X12 and X43) xor (X03 and X13 and X41) xor (X03 and X13 and X43) xor (X31 and X41) xor (X31 and X42) xor (X32 and X41) xor (X31 and X43) xor (X21 and X31 and X41) xor (X21 and X31 and X42) xor (X21 and X32 and X42) xor (X21 and X32 and X43) xor (X21 and X33 and X42) xor (X22 and X31 and X42) xor (X22 and X31 and X43) xor (X22 and X32 and X41) xor (X22 and X32 and X43) xor (X22 and X33 and X41) xor (X22 and X33 and X42) xor (X23 and X31 and X42) xor (X23 and X32 and X41) xor (X23 and X32 and X43) xor (X23 and X33 and X41) xor (X23 and X33 and X43) xor (X51) xor (X0_1 and X51) xor (X0_1 and X52) xor (X02 and X51) xor (X0_1 and X53) xor (X21 and X51) xor (X21 and X52) xor (X22 and X51) xor (X21 and X53) xor (X31 and X51) xor (X31 and X52) xor (X32 and X51) xor (X31 and X53) xor (X0_1 and X31 and X51) xor (X0_1 and X31 and X52) xor (X0_1 and X32 and X52) xor (X0_1 and X32 and X53) xor (X0_1 and X33 and X52) xor (X02 and X31 and X52) xor (X02 and X31 and X53) xor (X02 and X32 and X51) xor (X02 and X32 and X53) xor (X02 and X33 and X51) xor (X02 and X33 and X52) xor (X03 and X31 and X52) xor (X03 and X32 and X51) xor (X03 and X32 and X53) xor (X03 and X33 and X51) xor (X03 and X33 and X53) xor (X21 and X31 and X51) xor (X21 and X31 and X52) xor (X21 and X32 and X52) xor (X21 and X32 and X53) xor (X21 and X33 and X52) xor (X22 and X31 and X52) xor (X22 and X31 and X53) xor (X22 and X32 and X51) xor (X22 and X32 and X53) xor (X22 and X33 and X51) xor (X22 and X33 and X52) xor (X23 and X31 and X52) xor (X23 and X32 and X51) xor (X23 and X32 and X53) xor (X23 and X33 and X51) xor (X23 and X33 and X53) xor (X0_1 and X41 and X51) xor (X0_1 and X41 and X52) xor (X0_1 and X42 and X52) xor (X0_1 and X42 and X53) xor (X0_1 and X43 and X52) xor (X02 and X41 and X52) xor (X02 and X41 and X53) xor (X02 and X42 and X51) xor (X02 and X42 and X53) xor (X02 and X43 and X51) xor (X02 and X43 and X52) xor (X03 and X41 and X52) xor (X03 and X42 and X51) xor (X03 and X42 and X53) xor (X03 and X43 and X51) xor (X03 and X43 and X53) xor (X11 and X41 and X51) xor (X11 and X41 and X52) xor (X11 and X42 and X52) xor (X11 and X42 and X53) xor (X11 and X43 and X52) xor (X12 and X41 and X52) xor (X12 and X41 and X53) xor (X12 and X42 and X51) xor (X12 and X42 and X53) xor (X12 and X43 and X51) xor (X12 and X43 and X52) xor (X13 and X41 and X52) xor (X13 and X42 and X51) xor (X13 and X42 and X53) xor (X13 and X43 and X51) xor (X13 and X43 and X53) xor (X21 and X41 and X51) xor (X21 and X41 and X52) xor (X21 and X42 and X52) xor (X21 and X42 and X53) xor (X21 and X43 and X52) xor (X22 and X41 and X52) xor (X22 and X41 and X53) xor (X22 and X42 and X51) xor (X22 and X42 and X53) xor (X22 and X43 and X51) xor (X22 and X43 and X52) xor (X23 and X41 and X52) xor (X23 and X42 and X51) xor (X23 and X42 and X53) xor (X23 and X43 and X51) xor (X23 and X43 and X53) xor (X0_1 and X11 and X61) xor (X0_1 and X11 and X62) xor (X0_1 and X12 and X62) xor (X0_1 and X12 and X63) xor (X0_1 and X13 and X62) xor (X02 and X11 and X62) xor (X02 and X11 and X63) xor (X02 and X12 and X61) xor (X02 and X12 and X63) xor (X02 and X13 and X61) xor (X02 and X13 and X62) xor (X03 and X11 and X62) xor (X03 and X12 and X61) xor (X03 and X12 and X63) xor (X03 and X13 and X61) xor (X03 and X13 and X63) xor (X21 and X61) xor (X21 and X62) xor (X22 and X61) xor (X21 and X63) xor (X0_1 and X21 and X61) xor (X0_1 and X21 and X62) xor (X0_1 and X22 and X62) xor (X0_1 and X22 and X63) xor (X0_1 and X23 and X62) xor (X02 and X21 and X62) xor (X02 and X21 and X63) xor (X02 and X22 and X61) xor (X02 and X22 and X63) xor (X02 and X23 and X61) xor (X02 and X23 and X62) xor (X03 and X21 and X62) xor (X03 and X22 and X61) xor (X03 and X22 and X63) xor (X03 and X23 and X61) xor (X03 and X23 and X63) xor (X31 and X61) xor (X31 and X62) xor (X32 and X61) xor (X31 and X63) xor (X0_1 and X31 and X61) xor (X0_1 and X31 and X62) xor (X0_1 and X32 and X62) xor (X0_1 and X32 and X63) xor (X0_1 and X33 and X62) xor (X02 and X31 and X62) xor (X02 and X31 and X63) xor (X02 and X32 and X61) xor (X02 and X32 and X63) xor (X02 and X33 and X61) xor (X02 and X33 and X62) xor (X03 and X31 and X62) xor (X03 and X32 and X61) xor (X03 and X32 and X63) xor (X03 and X33 and X61) xor (X03 and X33 and X63) xor (X11 and X31 and X61) xor (X11 and X31 and X62) xor (X11 and X32 and X62) xor (X11 and X32 and X63) xor (X11 and X33 and X62) xor (X12 and X31 and X62) xor (X12 and X31 and X63) xor (X12 and X32 and X61) xor (X12 and X32 and X63) xor (X12 and X33 and X61) xor (X12 and X33 and X62) xor (X13 and X31 and X62) xor (X13 and X32 and X61) xor (X13 and X32 and X63) xor (X13 and X33 and X61) xor (X13 and X33 and X63) xor (X41 and X61) xor (X41 and X62) xor (X42 and X61) xor (X41 and X63) xor (X51 and X61) xor (X51 and X62) xor (X52 and X61) xor (X51 and X63) xor (X21 and X51 and X61) xor (X21 and X51 and X62) xor (X21 and X52 and X62) xor (X21 and X52 and X63) xor (X21 and X53 and X62) xor (X22 and X51 and X62) xor (X22 and X51 and X63) xor (X22 and X52 and X61) xor (X22 and X52 and X63) xor (X22 and X53 and X61) xor (X22 and X53 and X62) xor (X23 and X51 and X62) xor (X23 and X52 and X61) xor (X23 and X52 and X63) xor (X23 and X53 and X61) xor (X23 and X53 and X63) xor (X71) xor (X0_1 and X71) xor (X0_1 and X72) xor (X02 and X71) xor (X0_1 and X73) xor (X0_1 and X11 and X71) xor (X0_1 and X11 and X72) xor (X0_1 and X12 and X72) xor (X0_1 and X12 and X73) xor (X0_1 and X13 and X72) xor (X02 and X11 and X72) xor (X02 and X11 and X73) xor (X02 and X12 and X71) xor (X02 and X12 and X73) xor (X02 and X13 and X71) xor (X02 and X13 and X72) xor (X03 and X11 and X72) xor (X03 and X12 and X71) xor (X03 and X12 and X73) xor (X03 and X13 and X71) xor (X03 and X13 and X73) xor (X21 and X71) xor (X21 and X72) xor (X22 and X71) xor (X21 and X73) xor (X0_1 and X31 and X71) xor (X0_1 and X31 and X72) xor (X0_1 and X32 and X72) xor (X0_1 and X32 and X73) xor (X0_1 and X33 and X72) xor (X02 and X31 and X72) xor (X02 and X31 and X73) xor (X02 and X32 and X71) xor (X02 and X32 and X73) xor (X02 and X33 and X71) xor (X02 and X33 and X72) xor (X03 and X31 and X72) xor (X03 and X32 and X71) xor (X03 and X32 and X73) xor (X03 and X33 and X71) xor (X03 and X33 and X73) xor (X21 and X31 and X71) xor (X21 and X31 and X72) xor (X21 and X32 and X72) xor (X21 and X32 and X73) xor (X21 and X33 and X72) xor (X22 and X31 and X72) xor (X22 and X31 and X73) xor (X22 and X32 and X71) xor (X22 and X32 and X73) xor (X22 and X33 and X71) xor (X22 and X33 and X72) xor (X23 and X31 and X72) xor (X23 and X32 and X71) xor (X23 and X32 and X73) xor (X23 and X33 and X71) xor (X23 and X33 and X73) xor (X11 and X41 and X71) xor (X11 and X41 and X72) xor (X11 and X42 and X72) xor (X11 and X42 and X73) xor (X11 and X43 and X72) xor (X12 and X41 and X72) xor (X12 and X41 and X73) xor (X12 and X42 and X71) xor (X12 and X42 and X73) xor (X12 and X43 and X71) xor (X12 and X43 and X72) xor (X13 and X41 and X72) xor (X13 and X42 and X71) xor (X13 and X42 and X73) xor (X13 and X43 and X71) xor (X13 and X43 and X73) xor (X31 and X41 and X71) xor (X31 and X41 and X72) xor (X31 and X42 and X72) xor (X31 and X42 and X73) xor (X31 and X43 and X72) xor (X32 and X41 and X72) xor (X32 and X41 and X73) xor (X32 and X42 and X71) xor (X32 and X42 and X73) xor (X32 and X43 and X71) xor (X32 and X43 and X72) xor (X33 and X41 and X72) xor (X33 and X42 and X71) xor (X33 and X42 and X73) xor (X33 and X43 and X71) xor (X33 and X43 and X73) xor (X0_1 and X51 and X71) xor (X0_1 and X51 and X72) xor (X0_1 and X52 and X72) xor (X0_1 and X52 and X73) xor (X0_1 and X53 and X72) xor (X02 and X51 and X72) xor (X02 and X51 and X73) xor (X02 and X52 and X71) xor (X02 and X52 and X73) xor (X02 and X53 and X71) xor (X02 and X53 and X72) xor (X03 and X51 and X72) xor (X03 and X52 and X71) xor (X03 and X52 and X73) xor (X03 and X53 and X71) xor (X03 and X53 and X73) xor (X21 and X51 and X71) xor (X21 and X51 and X72) xor (X21 and X52 and X72) xor (X21 and X52 and X73) xor (X21 and X53 and X72) xor (X22 and X51 and X72) xor (X22 and X51 and X73) xor (X22 and X52 and X71) xor (X22 and X52 and X73) xor (X22 and X53 and X71) xor (X22 and X53 and X72) xor (X23 and X51 and X72) xor (X23 and X52 and X71) xor (X23 and X52 and X73) xor (X23 and X53 and X71) xor (X23 and X53 and X73) xor (X0_1 and X61 and X71) xor (X0_1 and X61 and X72) xor (X0_1 and X62 and X72) xor (X0_1 and X62 and X73) xor (X0_1 and X63 and X72) xor (X02 and X61 and X72) xor (X02 and X61 and X73) xor (X02 and X62 and X71) xor (X02 and X62 and X73) xor (X02 and X63 and X71) xor (X02 and X63 and X72) xor (X03 and X61 and X72) xor (X03 and X62 and X71) xor (X03 and X62 and X73) xor (X03 and X63 and X71) xor (X03 and X63 and X73) xor (X11 and X61 and X71) xor (X11 and X61 and X72) xor (X11 and X62 and X72) xor (X11 and X62 and X73) xor (X11 and X63 and X72) xor (X12 and X61 and X72) xor (X12 and X61 and X73) xor (X12 and X62 and X71) xor (X12 and X62 and X73) xor (X12 and X63 and X71) xor (X12 and X63 and X72) xor (X13 and X61 and X72) xor (X13 and X62 and X71) xor (X13 and X62 and X73) xor (X13 and X63 and X71) xor (X13 and X63 and X73) xor (X21 and X61 and X71) xor (X21 and X61 and X72) xor (X21 and X62 and X72) xor (X21 and X62 and X73) xor (X21 and X63 and X72) xor (X22 and X61 and X72) xor (X22 and X61 and X73) xor (X22 and X62 and X71) xor (X22 and X62 and X73) xor (X22 and X63 and X71) xor (X22 and X63 and X72) xor (X23 and X61 and X72) xor (X23 and X62 and X71) xor (X23 and X62 and X73) xor (X23 and X63 and X71) xor (X23 and X63 and X73) xor (X41 and X61 and X71) xor (X41 and X61 and X72) xor (X41 and X62 and X72) xor (X41 and X62 and X73) xor (X41 and X63 and X72) xor (X42 and X61 and X72) xor (X42 and X61 and X73) xor (X42 and X62 and X71) xor (X42 and X62 and X73) xor (X42 and X63 and X71) xor (X42 and X63 and X72) xor (X43 and X61 and X72) xor (X43 and X62 and X71) xor (X43 and X62 and X73) xor (X43 and X63 and X71) xor (X43 and X63 and X73));
    F02  <= ((X02) xor (X12) xor (X02 and X12) xor (X00 and X13) xor (X02 and X13) xor (X03 and X12) xor (X12 and X22) xor (X10 and X23) xor (X12 and X23) xor (X13 and X22) xor (X00 and X10 and X23) xor (X00 and X12 and X20) xor (X00 and X12 and X22) xor (X00 and X12 and X23) xor (X00 and X13 and X20) xor (X00 and X13 and X22) xor (X02 and X10 and X22) xor (X02 and X10 and X23) xor (X02 and X13 and X20) xor (X02 and X13 and X23) xor (X03 and X10 and X20) xor (X03 and X10 and X22) xor (X03 and X10 and X23) xor (X03 and X12 and X20) xor (X03 and X12 and X22) xor (X03 and X13 and X22) xor (X32) xor (X12 and X32) xor (X10 and X33) xor (X12 and X33) xor (X13 and X32) xor (X00 and X10 and X33) xor (X00 and X12 and X30) xor (X00 and X12 and X32) xor (X00 and X12 and X33) xor (X00 and X13 and X30) xor (X00 and X13 and X32) xor (X02 and X10 and X32) xor (X02 and X10 and X33) xor (X02 and X13 and X30) xor (X02 and X13 and X33) xor (X03 and X10 and X30) xor (X03 and X10 and X32) xor (X03 and X10 and X33) xor (X03 and X12 and X30) xor (X03 and X12 and X32) xor (X03 and X13 and X32) xor (X22 and X32) xor (X20 and X33) xor (X22 and X33) xor (X23 and X32) xor (X12 and X42) xor (X10 and X43) xor (X12 and X43) xor (X13 and X42) xor (X00 and X10 and X43) xor (X00 and X12 and X40) xor (X00 and X12 and X42) xor (X00 and X12 and X43) xor (X00 and X13 and X40) xor (X00 and X13 and X42) xor (X02 and X10 and X42) xor (X02 and X10 and X43) xor (X02 and X13 and X40) xor (X02 and X13 and X43) xor (X03 and X10 and X40) xor (X03 and X10 and X42) xor (X03 and X10 and X43) xor (X03 and X12 and X40) xor (X03 and X12 and X42) xor (X03 and X13 and X42) xor (X32 and X42) xor (X30 and X43) xor (X32 and X43) xor (X33 and X42) xor (X20 and X30 and X43) xor (X20 and X32 and X40) xor (X20 and X32 and X42) xor (X20 and X32 and X43) xor (X20 and X33 and X40) xor (X20 and X33 and X42) xor (X22 and X30 and X42) xor (X22 and X30 and X43) xor (X22 and X33 and X40) xor (X22 and X33 and X43) xor (X23 and X30 and X40) xor (X23 and X30 and X42) xor (X23 and X30 and X43) xor (X23 and X32 and X40) xor (X23 and X32 and X42) xor (X23 and X33 and X42) xor (X52) xor (X02 and X52) xor (X00 and X53) xor (X02 and X53) xor (X03 and X52) xor (X22 and X52) xor (X20 and X53) xor (X22 and X53) xor (X23 and X52) xor (X32 and X52) xor (X30 and X53) xor (X32 and X53) xor (X33 and X52) xor (X00 and X30 and X53) xor (X00 and X32 and X50) xor (X00 and X32 and X52) xor (X00 and X32 and X53) xor (X00 and X33 and X50) xor (X00 and X33 and X52) xor (X02 and X30 and X52) xor (X02 and X30 and X53) xor (X02 and X33 and X50) xor (X02 and X33 and X53) xor (X03 and X30 and X50) xor (X03 and X30 and X52) xor (X03 and X30 and X53) xor (X03 and X32 and X50) xor (X03 and X32 and X52) xor (X03 and X33 and X52) xor (X20 and X30 and X53) xor (X20 and X32 and X50) xor (X20 and X32 and X52) xor (X20 and X32 and X53) xor (X20 and X33 and X50) xor (X20 and X33 and X52) xor (X22 and X30 and X52) xor (X22 and X30 and X53) xor (X22 and X33 and X50) xor (X22 and X33 and X53) xor (X23 and X30 and X50) xor (X23 and X30 and X52) xor (X23 and X30 and X53) xor (X23 and X32 and X50) xor (X23 and X32 and X52) xor (X23 and X33 and X52) xor (X00 and X40 and X53) xor (X00 and X42 and X50) xor (X00 and X42 and X52) xor (X00 and X42 and X53) xor (X00 and X43 and X50) xor (X00 and X43 and X52) xor (X02 and X40 and X52) xor (X02 and X40 and X53) xor (X02 and X43 and X50) xor (X02 and X43 and X53) xor (X03 and X40 and X50) xor (X03 and X40 and X52) xor (X03 and X40 and X53) xor (X03 and X42 and X50) xor (X03 and X42 and X52) xor (X03 and X43 and X52) xor (X10 and X40 and X53) xor (X10 and X42 and X50) xor (X10 and X42 and X52) xor (X10 and X42 and X53) xor (X10 and X43 and X50) xor (X10 and X43 and X52) xor (X12 and X40 and X52) xor (X12 and X40 and X53) xor (X12 and X43 and X50) xor (X12 and X43 and X53) xor (X13 and X40 and X50) xor (X13 and X40 and X52) xor (X13 and X40 and X53) xor (X13 and X42 and X50) xor (X13 and X42 and X52) xor (X13 and X43 and X52) xor (X20 and X40 and X53) xor (X20 and X42 and X50) xor (X20 and X42 and X52) xor (X20 and X42 and X53) xor (X20 and X43 and X50) xor (X20 and X43 and X52) xor (X22 and X40 and X52) xor (X22 and X40 and X53) xor (X22 and X43 and X50) xor (X22 and X43 and X53) xor (X23 and X40 and X50) xor (X23 and X40 and X52) xor (X23 and X40 and X53) xor (X23 and X42 and X50) xor (X23 and X42 and X52) xor (X23 and X43 and X52) xor (X00 and X10 and X63) xor (X00 and X12 and X60) xor (X00 and X12 and X62) xor (X00 and X12 and X63) xor (X00 and X13 and X60) xor (X00 and X13 and X62) xor (X02 and X10 and X62) xor (X02 and X10 and X63) xor (X02 and X13 and X60) xor (X02 and X13 and X63) xor (X03 and X10 and X60) xor (X03 and X10 and X62) xor (X03 and X10 and X63) xor (X03 and X12 and X60) xor (X03 and X12 and X62) xor (X03 and X13 and X62) xor (X22 and X62) xor (X20 and X63) xor (X22 and X63) xor (X23 and X62) xor (X00 and X20 and X63) xor (X00 and X22 and X60) xor (X00 and X22 and X62) xor (X00 and X22 and X63) xor (X00 and X23 and X60) xor (X00 and X23 and X62) xor (X02 and X20 and X62) xor (X02 and X20 and X63) xor (X02 and X23 and X60) xor (X02 and X23 and X63) xor (X03 and X20 and X60) xor (X03 and X20 and X62) xor (X03 and X20 and X63) xor (X03 and X22 and X60) xor (X03 and X22 and X62) xor (X03 and X23 and X62) xor (X32 and X62) xor (X30 and X63) xor (X32 and X63) xor (X33 and X62) xor (X00 and X30 and X63) xor (X00 and X32 and X60) xor (X00 and X32 and X62) xor (X00 and X32 and X63) xor (X00 and X33 and X60) xor (X00 and X33 and X62) xor (X02 and X30 and X62) xor (X02 and X30 and X63) xor (X02 and X33 and X60) xor (X02 and X33 and X63) xor (X03 and X30 and X60) xor (X03 and X30 and X62) xor (X03 and X30 and X63) xor (X03 and X32 and X60) xor (X03 and X32 and X62) xor (X03 and X33 and X62) xor (X10 and X30 and X63) xor (X10 and X32 and X60) xor (X10 and X32 and X62) xor (X10 and X32 and X63) xor (X10 and X33 and X60) xor (X10 and X33 and X62) xor (X12 and X30 and X62) xor (X12 and X30 and X63) xor (X12 and X33 and X60) xor (X12 and X33 and X63) xor (X13 and X30 and X60) xor (X13 and X30 and X62) xor (X13 and X30 and X63) xor (X13 and X32 and X60) xor (X13 and X32 and X62) xor (X13 and X33 and X62) xor (X42 and X62) xor (X40 and X63) xor (X42 and X63) xor (X43 and X62) xor (X52 and X62) xor (X50 and X63) xor (X52 and X63) xor (X53 and X62) xor (X20 and X50 and X63) xor (X20 and X52 and X60) xor (X20 and X52 and X62) xor (X20 and X52 and X63) xor (X20 and X53 and X60) xor (X20 and X53 and X62) xor (X22 and X50 and X62) xor (X22 and X50 and X63) xor (X22 and X53 and X60) xor (X22 and X53 and X63) xor (X23 and X50 and X60) xor (X23 and X50 and X62) xor (X23 and X50 and X63) xor (X23 and X52 and X60) xor (X23 and X52 and X62) xor (X23 and X53 and X62) xor (X72) xor (X02 and X72) xor (X00 and X73) xor (X02 and X73) xor (X03 and X72) xor (X00 and X10 and X73) xor (X00 and X12 and X70) xor (X00 and X12 and X72) xor (X00 and X12 and X73) xor (X00 and X13 and X70) xor (X00 and X13 and X72) xor (X02 and X10 and X72) xor (X02 and X10 and X73) xor (X02 and X13 and X70) xor (X02 and X13 and X73) xor (X03 and X10 and X70) xor (X03 and X10 and X72) xor (X03 and X10 and X73) xor (X03 and X12 and X70) xor (X03 and X12 and X72) xor (X03 and X13 and X72) xor (X22 and X72) xor (X20 and X73) xor (X22 and X73) xor (X23 and X72) xor (X00 and X30 and X73) xor (X00 and X32 and X70) xor (X00 and X32 and X72) xor (X00 and X32 and X73) xor (X00 and X33 and X70) xor (X00 and X33 and X72) xor (X02 and X30 and X72) xor (X02 and X30 and X73) xor (X02 and X33 and X70) xor (X02 and X33 and X73) xor (X03 and X30 and X70) xor (X03 and X30 and X72) xor (X03 and X30 and X73) xor (X03 and X32 and X70) xor (X03 and X32 and X72) xor (X03 and X33 and X72) xor (X20 and X30 and X73) xor (X20 and X32 and X70) xor (X20 and X32 and X72) xor (X20 and X32 and X73) xor (X20 and X33 and X70) xor (X20 and X33 and X72) xor (X22 and X30 and X72) xor (X22 and X30 and X73) xor (X22 and X33 and X70) xor (X22 and X33 and X73) xor (X23 and X30 and X70) xor (X23 and X30 and X72) xor (X23 and X30 and X73) xor (X23 and X32 and X70) xor (X23 and X32 and X72) xor (X23 and X33 and X72) xor (X10 and X40 and X73) xor (X10 and X42 and X70) xor (X10 and X42 and X72) xor (X10 and X42 and X73) xor (X10 and X43 and X70) xor (X10 and X43 and X72) xor (X12 and X40 and X72) xor (X12 and X40 and X73) xor (X12 and X43 and X70) xor (X12 and X43 and X73) xor (X13 and X40 and X70) xor (X13 and X40 and X72) xor (X13 and X40 and X73) xor (X13 and X42 and X70) xor (X13 and X42 and X72) xor (X13 and X43 and X72) xor (X30 and X40 and X73) xor (X30 and X42 and X70) xor (X30 and X42 and X72) xor (X30 and X42 and X73) xor (X30 and X43 and X70) xor (X30 and X43 and X72) xor (X32 and X40 and X72) xor (X32 and X40 and X73) xor (X32 and X43 and X70) xor (X32 and X43 and X73) xor (X33 and X40 and X70) xor (X33 and X40 and X72) xor (X33 and X40 and X73) xor (X33 and X42 and X70) xor (X33 and X42 and X72) xor (X33 and X43 and X72) xor (X00 and X50 and X73) xor (X00 and X52 and X70) xor (X00 and X52 and X72) xor (X00 and X52 and X73) xor (X00 and X53 and X70) xor (X00 and X53 and X72) xor (X02 and X50 and X72) xor (X02 and X50 and X73) xor (X02 and X53 and X70) xor (X02 and X53 and X73) xor (X03 and X50 and X70) xor (X03 and X50 and X72) xor (X03 and X50 and X73) xor (X03 and X52 and X70) xor (X03 and X52 and X72) xor (X03 and X53 and X72) xor (X20 and X50 and X73) xor (X20 and X52 and X70) xor (X20 and X52 and X72) xor (X20 and X52 and X73) xor (X20 and X53 and X70) xor (X20 and X53 and X72) xor (X22 and X50 and X72) xor (X22 and X50 and X73) xor (X22 and X53 and X70) xor (X22 and X53 and X73) xor (X23 and X50 and X70) xor (X23 and X50 and X72) xor (X23 and X50 and X73) xor (X23 and X52 and X70) xor (X23 and X52 and X72) xor (X23 and X53 and X72) xor (X00 and X60 and X73) xor (X00 and X62 and X70) xor (X00 and X62 and X72) xor (X00 and X62 and X73) xor (X00 and X63 and X70) xor (X00 and X63 and X72) xor (X02 and X60 and X72) xor (X02 and X60 and X73) xor (X02 and X63 and X70) xor (X02 and X63 and X73) xor (X03 and X60 and X70) xor (X03 and X60 and X72) xor (X03 and X60 and X73) xor (X03 and X62 and X70) xor (X03 and X62 and X72) xor (X03 and X63 and X72) xor (X10 and X60 and X73) xor (X10 and X62 and X70) xor (X10 and X62 and X72) xor (X10 and X62 and X73) xor (X10 and X63 and X70) xor (X10 and X63 and X72) xor (X12 and X60 and X72) xor (X12 and X60 and X73) xor (X12 and X63 and X70) xor (X12 and X63 and X73) xor (X13 and X60 and X70) xor (X13 and X60 and X72) xor (X13 and X60 and X73) xor (X13 and X62 and X70) xor (X13 and X62 and X72) xor (X13 and X63 and X72) xor (X20 and X60 and X73) xor (X20 and X62 and X70) xor (X20 and X62 and X72) xor (X20 and X62 and X73) xor (X20 and X63 and X70) xor (X20 and X63 and X72) xor (X22 and X60 and X72) xor (X22 and X60 and X73) xor (X22 and X63 and X70) xor (X22 and X63 and X73) xor (X23 and X60 and X70) xor (X23 and X60 and X72) xor (X23 and X60 and X73) xor (X23 and X62 and X70) xor (X23 and X62 and X72) xor (X23 and X63 and X72) xor (X40 and X60 and X73) xor (X40 and X62 and X70) xor (X40 and X62 and X72) xor (X40 and X62 and X73) xor (X40 and X63 and X70) xor (X40 and X63 and X72) xor (X42 and X60 and X72) xor (X42 and X60 and X73) xor (X42 and X63 and X70) xor (X42 and X63 and X73) xor (X43 and X60 and X70) xor (X43 and X60 and X72) xor (X43 and X60 and X73) xor (X43 and X62 and X70) xor (X43 and X62 and X72) xor (X43 and X63 and X72));
    F03  <= ((X03) xor (X13) xor (X03 and X13) xor (X03 and X10) xor (X03 and X11) xor (X0_1 and X10) xor (X13 and X23) xor (X13 and X20) xor (X13 and X21) xor (X11 and X20) xor (X00 and X10 and X21) xor (X00 and X11 and X20) xor (X00 and X11 and X23) xor (X00 and X13 and X21) xor (X00 and X13 and X23) xor (X0_1 and X10 and X21) xor (X0_1 and X10 and X23) xor (X0_1 and X11 and X23) xor (X0_1 and X13 and X20) xor (X0_1 and X13 and X21) xor (X0_1 and X13 and X23) xor (X03 and X10 and X21) xor (X03 and X11 and X20) xor (X03 and X11 and X21) xor (X03 and X11 and X23) xor (X03 and X13 and X20) xor (X33) xor (X13 and X33) xor (X13 and X30) xor (X13 and X31) xor (X11 and X30) xor (X00 and X10 and X31) xor (X00 and X11 and X30) xor (X00 and X11 and X33) xor (X00 and X13 and X31) xor (X00 and X13 and X33) xor (X0_1 and X10 and X31) xor (X0_1 and X10 and X33) xor (X0_1 and X11 and X33) xor (X0_1 and X13 and X30) xor (X0_1 and X13 and X31) xor (X0_1 and X13 and X33) xor (X03 and X10 and X31) xor (X03 and X11 and X30) xor (X03 and X11 and X31) xor (X03 and X11 and X33) xor (X03 and X13 and X30) xor (X23 and X33) xor (X23 and X30) xor (X23 and X31) xor (X21 and X30) xor (X13 and X43) xor (X13 and X40) xor (X13 and X41) xor (X11 and X40) xor (X00 and X10 and X41) xor (X00 and X11 and X40) xor (X00 and X11 and X43) xor (X00 and X13 and X41) xor (X00 and X13 and X43) xor (X0_1 and X10 and X41) xor (X0_1 and X10 and X43) xor (X0_1 and X11 and X43) xor (X0_1 and X13 and X40) xor (X0_1 and X13 and X41) xor (X0_1 and X13 and X43) xor (X03 and X10 and X41) xor (X03 and X11 and X40) xor (X03 and X11 and X41) xor (X03 and X11 and X43) xor (X03 and X13 and X40) xor (X33 and X43) xor (X33 and X40) xor (X33 and X41) xor (X31 and X40) xor (X20 and X30 and X41) xor (X20 and X31 and X40) xor (X20 and X31 and X43) xor (X20 and X33 and X41) xor (X20 and X33 and X43) xor (X21 and X30 and X41) xor (X21 and X30 and X43) xor (X21 and X31 and X43) xor (X21 and X33 and X40) xor (X21 and X33 and X41) xor (X21 and X33 and X43) xor (X23 and X30 and X41) xor (X23 and X31 and X40) xor (X23 and X31 and X41) xor (X23 and X31 and X43) xor (X23 and X33 and X40) xor (X53) xor (X03 and X53) xor (X03 and X50) xor (X03 and X51) xor (X0_1 and X50) xor (X23 and X53) xor (X23 and X50) xor (X23 and X51) xor (X21 and X50) xor (X33 and X53) xor (X33 and X50) xor (X33 and X51) xor (X31 and X50) xor (X00 and X30 and X51) xor (X00 and X31 and X50) xor (X00 and X31 and X53) xor (X00 and X33 and X51) xor (X00 and X33 and X53) xor (X0_1 and X30 and X51) xor (X0_1 and X30 and X53) xor (X0_1 and X31 and X53) xor (X0_1 and X33 and X50) xor (X0_1 and X33 and X51) xor (X0_1 and X33 and X53) xor (X03 and X30 and X51) xor (X03 and X31 and X50) xor (X03 and X31 and X51) xor (X03 and X31 and X53) xor (X03 and X33 and X50) xor (X20 and X30 and X51) xor (X20 and X31 and X50) xor (X20 and X31 and X53) xor (X20 and X33 and X51) xor (X20 and X33 and X53) xor (X21 and X30 and X51) xor (X21 and X30 and X53) xor (X21 and X31 and X53) xor (X21 and X33 and X50) xor (X21 and X33 and X51) xor (X21 and X33 and X53) xor (X23 and X30 and X51) xor (X23 and X31 and X50) xor (X23 and X31 and X51) xor (X23 and X31 and X53) xor (X23 and X33 and X50) xor (X00 and X40 and X51) xor (X00 and X41 and X50) xor (X00 and X41 and X53) xor (X00 and X43 and X51) xor (X00 and X43 and X53) xor (X0_1 and X40 and X51) xor (X0_1 and X40 and X53) xor (X0_1 and X41 and X53) xor (X0_1 and X43 and X50) xor (X0_1 and X43 and X51) xor (X0_1 and X43 and X53) xor (X03 and X40 and X51) xor (X03 and X41 and X50) xor (X03 and X41 and X51) xor (X03 and X41 and X53) xor (X03 and X43 and X50) xor (X10 and X40 and X51) xor (X10 and X41 and X50) xor (X10 and X41 and X53) xor (X10 and X43 and X51) xor (X10 and X43 and X53) xor (X11 and X40 and X51) xor (X11 and X40 and X53) xor (X11 and X41 and X53) xor (X11 and X43 and X50) xor (X11 and X43 and X51) xor (X11 and X43 and X53) xor (X13 and X40 and X51) xor (X13 and X41 and X50) xor (X13 and X41 and X51) xor (X13 and X41 and X53) xor (X13 and X43 and X50) xor (X20 and X40 and X51) xor (X20 and X41 and X50) xor (X20 and X41 and X53) xor (X20 and X43 and X51) xor (X20 and X43 and X53) xor (X21 and X40 and X51) xor (X21 and X40 and X53) xor (X21 and X41 and X53) xor (X21 and X43 and X50) xor (X21 and X43 and X51) xor (X21 and X43 and X53) xor (X23 and X40 and X51) xor (X23 and X41 and X50) xor (X23 and X41 and X51) xor (X23 and X41 and X53) xor (X23 and X43 and X50) xor (X00 and X10 and X61) xor (X00 and X11 and X60) xor (X00 and X11 and X63) xor (X00 and X13 and X61) xor (X00 and X13 and X63) xor (X0_1 and X10 and X61) xor (X0_1 and X10 and X63) xor (X0_1 and X11 and X63) xor (X0_1 and X13 and X60) xor (X0_1 and X13 and X61) xor (X0_1 and X13 and X63) xor (X03 and X10 and X61) xor (X03 and X11 and X60) xor (X03 and X11 and X61) xor (X03 and X11 and X63) xor (X03 and X13 and X60) xor (X23 and X63) xor (X23 and X60) xor (X23 and X61) xor (X21 and X60) xor (X00 and X20 and X61) xor (X00 and X21 and X60) xor (X00 and X21 and X63) xor (X00 and X23 and X61) xor (X00 and X23 and X63) xor (X0_1 and X20 and X61) xor (X0_1 and X20 and X63) xor (X0_1 and X21 and X63) xor (X0_1 and X23 and X60) xor (X0_1 and X23 and X61) xor (X0_1 and X23 and X63) xor (X03 and X20 and X61) xor (X03 and X21 and X60) xor (X03 and X21 and X61) xor (X03 and X21 and X63) xor (X03 and X23 and X60) xor (X33 and X63) xor (X33 and X60) xor (X33 and X61) xor (X31 and X60) xor (X00 and X30 and X61) xor (X00 and X31 and X60) xor (X00 and X31 and X63) xor (X00 and X33 and X61) xor (X00 and X33 and X63) xor (X0_1 and X30 and X61) xor (X0_1 and X30 and X63) xor (X0_1 and X31 and X63) xor (X0_1 and X33 and X60) xor (X0_1 and X33 and X61) xor (X0_1 and X33 and X63) xor (X03 and X30 and X61) xor (X03 and X31 and X60) xor (X03 and X31 and X61) xor (X03 and X31 and X63) xor (X03 and X33 and X60) xor (X10 and X30 and X61) xor (X10 and X31 and X60) xor (X10 and X31 and X63) xor (X10 and X33 and X61) xor (X10 and X33 and X63) xor (X11 and X30 and X61) xor (X11 and X30 and X63) xor (X11 and X31 and X63) xor (X11 and X33 and X60) xor (X11 and X33 and X61) xor (X11 and X33 and X63) xor (X13 and X30 and X61) xor (X13 and X31 and X60) xor (X13 and X31 and X61) xor (X13 and X31 and X63) xor (X13 and X33 and X60) xor (X43 and X63) xor (X43 and X60) xor (X43 and X61) xor (X41 and X60) xor (X53 and X63) xor (X53 and X60) xor (X53 and X61) xor (X51 and X60) xor (X20 and X50 and X61) xor (X20 and X51 and X60) xor (X20 and X51 and X63) xor (X20 and X53 and X61) xor (X20 and X53 and X63) xor (X21 and X50 and X61) xor (X21 and X50 and X63) xor (X21 and X51 and X63) xor (X21 and X53 and X60) xor (X21 and X53 and X61) xor (X21 and X53 and X63) xor (X23 and X50 and X61) xor (X23 and X51 and X60) xor (X23 and X51 and X61) xor (X23 and X51 and X63) xor (X23 and X53 and X60) xor (X73) xor (X03 and X73) xor (X03 and X70) xor (X03 and X71) xor (X0_1 and X70) xor (X00 and X10 and X71) xor (X00 and X11 and X70) xor (X00 and X11 and X73) xor (X00 and X13 and X71) xor (X00 and X13 and X73) xor (X0_1 and X10 and X71) xor (X0_1 and X10 and X73) xor (X0_1 and X11 and X73) xor (X0_1 and X13 and X70) xor (X0_1 and X13 and X71) xor (X0_1 and X13 and X73) xor (X03 and X10 and X71) xor (X03 and X11 and X70) xor (X03 and X11 and X71) xor (X03 and X11 and X73) xor (X03 and X13 and X70) xor (X23 and X73) xor (X23 and X70) xor (X23 and X71) xor (X21 and X70) xor (X00 and X30 and X71) xor (X00 and X31 and X70) xor (X00 and X31 and X73) xor (X00 and X33 and X71) xor (X00 and X33 and X73) xor (X0_1 and X30 and X71) xor (X0_1 and X30 and X73) xor (X0_1 and X31 and X73) xor (X0_1 and X33 and X70) xor (X0_1 and X33 and X71) xor (X0_1 and X33 and X73) xor (X03 and X30 and X71) xor (X03 and X31 and X70) xor (X03 and X31 and X71) xor (X03 and X31 and X73) xor (X03 and X33 and X70) xor (X20 and X30 and X71) xor (X20 and X31 and X70) xor (X20 and X31 and X73) xor (X20 and X33 and X71) xor (X20 and X33 and X73) xor (X21 and X30 and X71) xor (X21 and X30 and X73) xor (X21 and X31 and X73) xor (X21 and X33 and X70) xor (X21 and X33 and X71) xor (X21 and X33 and X73) xor (X23 and X30 and X71) xor (X23 and X31 and X70) xor (X23 and X31 and X71) xor (X23 and X31 and X73) xor (X23 and X33 and X70) xor (X10 and X40 and X71) xor (X10 and X41 and X70) xor (X10 and X41 and X73) xor (X10 and X43 and X71) xor (X10 and X43 and X73) xor (X11 and X40 and X71) xor (X11 and X40 and X73) xor (X11 and X41 and X73) xor (X11 and X43 and X70) xor (X11 and X43 and X71) xor (X11 and X43 and X73) xor (X13 and X40 and X71) xor (X13 and X41 and X70) xor (X13 and X41 and X71) xor (X13 and X41 and X73) xor (X13 and X43 and X70) xor (X30 and X40 and X71) xor (X30 and X41 and X70) xor (X30 and X41 and X73) xor (X30 and X43 and X71) xor (X30 and X43 and X73) xor (X31 and X40 and X71) xor (X31 and X40 and X73) xor (X31 and X41 and X73) xor (X31 and X43 and X70) xor (X31 and X43 and X71) xor (X31 and X43 and X73) xor (X33 and X40 and X71) xor (X33 and X41 and X70) xor (X33 and X41 and X71) xor (X33 and X41 and X73) xor (X33 and X43 and X70) xor (X00 and X50 and X71) xor (X00 and X51 and X70) xor (X00 and X51 and X73) xor (X00 and X53 and X71) xor (X00 and X53 and X73) xor (X0_1 and X50 and X71) xor (X0_1 and X50 and X73) xor (X0_1 and X51 and X73) xor (X0_1 and X53 and X70) xor (X0_1 and X53 and X71) xor (X0_1 and X53 and X73) xor (X03 and X50 and X71) xor (X03 and X51 and X70) xor (X03 and X51 and X71) xor (X03 and X51 and X73) xor (X03 and X53 and X70) xor (X20 and X50 and X71) xor (X20 and X51 and X70) xor (X20 and X51 and X73) xor (X20 and X53 and X71) xor (X20 and X53 and X73) xor (X21 and X50 and X71) xor (X21 and X50 and X73) xor (X21 and X51 and X73) xor (X21 and X53 and X70) xor (X21 and X53 and X71) xor (X21 and X53 and X73) xor (X23 and X50 and X71) xor (X23 and X51 and X70) xor (X23 and X51 and X71) xor (X23 and X51 and X73) xor (X23 and X53 and X70) xor (X00 and X60 and X71) xor (X00 and X61 and X70) xor (X00 and X61 and X73) xor (X00 and X63 and X71) xor (X00 and X63 and X73) xor (X0_1 and X60 and X71) xor (X0_1 and X60 and X73) xor (X0_1 and X61 and X73) xor (X0_1 and X63 and X70) xor (X0_1 and X63 and X71) xor (X0_1 and X63 and X73) xor (X03 and X60 and X71) xor (X03 and X61 and X70) xor (X03 and X61 and X71) xor (X03 and X61 and X73) xor (X03 and X63 and X70) xor (X10 and X60 and X71) xor (X10 and X61 and X70) xor (X10 and X61 and X73) xor (X10 and X63 and X71) xor (X10 and X63 and X73) xor (X11 and X60 and X71) xor (X11 and X60 and X73) xor (X11 and X61 and X73) xor (X11 and X63 and X70) xor (X11 and X63 and X71) xor (X11 and X63 and X73) xor (X13 and X60 and X71) xor (X13 and X61 and X70) xor (X13 and X61 and X71) xor (X13 and X61 and X73) xor (X13 and X63 and X70) xor (X20 and X60 and X71) xor (X20 and X61 and X70) xor (X20 and X61 and X73) xor (X20 and X63 and X71) xor (X20 and X63 and X73) xor (X21 and X60 and X71) xor (X21 and X60 and X73) xor (X21 and X61 and X73) xor (X21 and X63 and X70) xor (X21 and X63 and X71) xor (X21 and X63 and X73) xor (X23 and X60 and X71) xor (X23 and X61 and X70) xor (X23 and X61 and X71) xor (X23 and X61 and X73) xor (X23 and X63 and X70) xor (X40 and X60 and X71) xor (X40 and X61 and X70) xor (X40 and X61 and X73) xor (X40 and X63 and X71) xor (X40 and X63 and X73) xor (X41 and X60 and X71) xor (X41 and X60 and X73) xor (X41 and X61 and X73) xor (X41 and X63 and X70) xor (X41 and X63 and X71) xor (X41 and X63 and X73) xor (X43 and X60 and X71) xor (X43 and X61 and X70) xor (X43 and X61 and X71) xor (X43 and X61 and X73) xor (X43 and X63 and X70));
    F10  <= ((X10) xor (X00 and X10) xor (X00 and X11) xor (X02 and X10) xor (X00 and X12) xor (X00 and X20) xor (X00 and X21) xor (X02 and X20) xor (X00 and X22) xor (X00 and X10 and X20) xor (X00 and X10 and X22) xor (X00 and X11 and X21) xor (X00 and X11 and X22) xor (X00 and X12 and X21) xor (X0_1 and X10 and X20) xor (X0_1 and X10 and X22) xor (X0_1 and X11 and X20) xor (X0_1 and X12 and X20) xor (X0_1 and X12 and X21) xor (X02 and X10 and X20) xor (X02 and X10 and X21) xor (X02 and X11 and X20) xor (X02 and X11 and X21) xor (X02 and X12 and X20) xor (X02 and X12 and X22) xor (X00 and X30) xor (X00 and X31) xor (X02 and X30) xor (X00 and X32) xor (X00 and X10 and X30) xor (X00 and X10 and X32) xor (X00 and X11 and X31) xor (X00 and X11 and X32) xor (X00 and X12 and X31) xor (X0_1 and X10 and X30) xor (X0_1 and X10 and X32) xor (X0_1 and X11 and X30) xor (X0_1 and X12 and X30) xor (X0_1 and X12 and X31) xor (X02 and X10 and X30) xor (X02 and X10 and X31) xor (X02 and X11 and X30) xor (X02 and X11 and X31) xor (X02 and X12 and X30) xor (X02 and X12 and X32) xor (X00 and X10 and X40) xor (X00 and X10 and X42) xor (X00 and X11 and X41) xor (X00 and X11 and X42) xor (X00 and X12 and X41) xor (X0_1 and X10 and X40) xor (X0_1 and X10 and X42) xor (X0_1 and X11 and X40) xor (X0_1 and X12 and X40) xor (X0_1 and X12 and X41) xor (X02 and X10 and X40) xor (X02 and X10 and X41) xor (X02 and X11 and X40) xor (X02 and X11 and X41) xor (X02 and X12 and X40) xor (X02 and X12 and X42) xor (X20 and X40) xor (X20 and X41) xor (X22 and X40) xor (X20 and X42) xor (X00 and X20 and X40) xor (X00 and X20 and X42) xor (X00 and X21 and X41) xor (X00 and X21 and X42) xor (X00 and X22 and X41) xor (X0_1 and X20 and X40) xor (X0_1 and X20 and X42) xor (X0_1 and X21 and X40) xor (X0_1 and X22 and X40) xor (X0_1 and X22 and X41) xor (X02 and X20 and X40) xor (X02 and X20 and X41) xor (X02 and X21 and X40) xor (X02 and X21 and X41) xor (X02 and X22 and X40) xor (X02 and X22 and X42) xor (X00 and X30 and X40) xor (X00 and X30 and X42) xor (X00 and X31 and X41) xor (X00 and X31 and X42) xor (X00 and X32 and X41) xor (X0_1 and X30 and X40) xor (X0_1 and X30 and X42) xor (X0_1 and X31 and X40) xor (X0_1 and X32 and X40) xor (X0_1 and X32 and X41) xor (X02 and X30 and X40) xor (X02 and X30 and X41) xor (X02 and X31 and X40) xor (X02 and X31 and X41) xor (X02 and X32 and X40) xor (X02 and X32 and X42) xor (X50) xor (X10 and X50) xor (X10 and X51) xor (X12 and X50) xor (X10 and X52) xor (X20 and X50) xor (X20 and X51) xor (X22 and X50) xor (X20 and X52) xor (X30 and X50) xor (X30 and X51) xor (X32 and X50) xor (X30 and X52) xor (X10 and X30 and X50) xor (X10 and X30 and X52) xor (X10 and X31 and X51) xor (X10 and X31 and X52) xor (X10 and X32 and X51) xor (X11 and X30 and X50) xor (X11 and X30 and X52) xor (X11 and X31 and X50) xor (X11 and X32 and X50) xor (X11 and X32 and X51) xor (X12 and X30 and X50) xor (X12 and X30 and X51) xor (X12 and X31 and X50) xor (X12 and X31 and X51) xor (X12 and X32 and X50) xor (X12 and X32 and X52) xor (X20 and X30 and X50) xor (X20 and X30 and X52) xor (X20 and X31 and X51) xor (X20 and X31 and X52) xor (X20 and X32 and X51) xor (X21 and X30 and X50) xor (X21 and X30 and X52) xor (X21 and X31 and X50) xor (X21 and X32 and X50) xor (X21 and X32 and X51) xor (X22 and X30 and X50) xor (X22 and X30 and X51) xor (X22 and X31 and X50) xor (X22 and X31 and X51) xor (X22 and X32 and X50) xor (X22 and X32 and X52) xor (X30 and X40 and X50) xor (X30 and X40 and X52) xor (X30 and X41 and X51) xor (X30 and X41 and X52) xor (X30 and X42 and X51) xor (X31 and X40 and X50) xor (X31 and X40 and X52) xor (X31 and X41 and X50) xor (X31 and X42 and X50) xor (X31 and X42 and X51) xor (X32 and X40 and X50) xor (X32 and X40 and X51) xor (X32 and X41 and X50) xor (X32 and X41 and X51) xor (X32 and X42 and X50) xor (X32 and X42 and X52) xor (X60) xor (X10 and X60) xor (X10 and X61) xor (X12 and X60) xor (X10 and X62) xor (X00 and X10 and X60) xor (X00 and X10 and X62) xor (X00 and X11 and X61) xor (X00 and X11 and X62) xor (X00 and X12 and X61) xor (X0_1 and X10 and X60) xor (X0_1 and X10 and X62) xor (X0_1 and X11 and X60) xor (X0_1 and X12 and X60) xor (X0_1 and X12 and X61) xor (X02 and X10 and X60) xor (X02 and X10 and X61) xor (X02 and X11 and X60) xor (X02 and X11 and X61) xor (X02 and X12 and X60) xor (X02 and X12 and X62) xor (X20 and X60) xor (X20 and X61) xor (X22 and X60) xor (X20 and X62) xor (X00 and X20 and X60) xor (X00 and X20 and X62) xor (X00 and X21 and X61) xor (X00 and X21 and X62) xor (X00 and X22 and X61) xor (X0_1 and X20 and X60) xor (X0_1 and X20 and X62) xor (X0_1 and X21 and X60) xor (X0_1 and X22 and X60) xor (X0_1 and X22 and X61) xor (X02 and X20 and X60) xor (X02 and X20 and X61) xor (X02 and X21 and X60) xor (X02 and X21 and X61) xor (X02 and X22 and X60) xor (X02 and X22 and X62) xor (X00 and X30 and X60) xor (X00 and X30 and X62) xor (X00 and X31 and X61) xor (X00 and X31 and X62) xor (X00 and X32 and X61) xor (X0_1 and X30 and X60) xor (X0_1 and X30 and X62) xor (X0_1 and X31 and X60) xor (X0_1 and X32 and X60) xor (X0_1 and X32 and X61) xor (X02 and X30 and X60) xor (X02 and X30 and X61) xor (X02 and X31 and X60) xor (X02 and X31 and X61) xor (X02 and X32 and X60) xor (X02 and X32 and X62) xor (X40 and X60) xor (X40 and X61) xor (X42 and X60) xor (X40 and X62) xor (X10 and X40 and X60) xor (X10 and X40 and X62) xor (X10 and X41 and X61) xor (X10 and X41 and X62) xor (X10 and X42 and X61) xor (X11 and X40 and X60) xor (X11 and X40 and X62) xor (X11 and X41 and X60) xor (X11 and X42 and X60) xor (X11 and X42 and X61) xor (X12 and X40 and X60) xor (X12 and X40 and X61) xor (X12 and X41 and X60) xor (X12 and X41 and X61) xor (X12 and X42 and X60) xor (X12 and X42 and X62) xor (X30 and X50 and X60) xor (X30 and X50 and X62) xor (X30 and X51 and X61) xor (X30 and X51 and X62) xor (X30 and X52 and X61) xor (X31 and X50 and X60) xor (X31 and X50 and X62) xor (X31 and X51 and X60) xor (X31 and X52 and X60) xor (X31 and X52 and X61) xor (X32 and X50 and X60) xor (X32 and X50 and X61) xor (X32 and X51 and X60) xor (X32 and X51 and X61) xor (X32 and X52 and X60) xor (X32 and X52 and X62) xor (X40 and X50 and X60) xor (X40 and X50 and X62) xor (X40 and X51 and X61) xor (X40 and X51 and X62) xor (X40 and X52 and X61) xor (X41 and X50 and X60) xor (X41 and X50 and X62) xor (X41 and X51 and X60) xor (X41 and X52 and X60) xor (X41 and X52 and X61) xor (X42 and X50 and X60) xor (X42 and X50 and X61) xor (X42 and X51 and X60) xor (X42 and X51 and X61) xor (X42 and X52 and X60) xor (X42 and X52 and X62) xor (X70) xor (X10 and X70) xor (X10 and X71) xor (X12 and X70) xor (X10 and X72) xor (X00 and X10 and X70) xor (X00 and X10 and X72) xor (X00 and X11 and X71) xor (X00 and X11 and X72) xor (X00 and X12 and X71) xor (X0_1 and X10 and X70) xor (X0_1 and X10 and X72) xor (X0_1 and X11 and X70) xor (X0_1 and X12 and X70) xor (X0_1 and X12 and X71) xor (X02 and X10 and X70) xor (X02 and X10 and X71) xor (X02 and X11 and X70) xor (X02 and X11 and X71) xor (X02 and X12 and X70) xor (X02 and X12 and X72) xor (X00 and X20 and X70) xor (X00 and X20 and X72) xor (X00 and X21 and X71) xor (X00 and X21 and X72) xor (X00 and X22 and X71) xor (X0_1 and X20 and X70) xor (X0_1 and X20 and X72) xor (X0_1 and X21 and X70) xor (X0_1 and X22 and X70) xor (X0_1 and X22 and X71) xor (X02 and X20 and X70) xor (X02 and X20 and X71) xor (X02 and X21 and X70) xor (X02 and X21 and X71) xor (X02 and X22 and X70) xor (X02 and X22 and X72) xor (X00 and X30 and X70) xor (X00 and X30 and X72) xor (X00 and X31 and X71) xor (X00 and X31 and X72) xor (X00 and X32 and X71) xor (X0_1 and X30 and X70) xor (X0_1 and X30 and X72) xor (X0_1 and X31 and X70) xor (X0_1 and X32 and X70) xor (X0_1 and X32 and X71) xor (X02 and X30 and X70) xor (X02 and X30 and X71) xor (X02 and X31 and X70) xor (X02 and X31 and X71) xor (X02 and X32 and X70) xor (X02 and X32 and X72) xor (X10 and X30 and X70) xor (X10 and X30 and X72) xor (X10 and X31 and X71) xor (X10 and X31 and X72) xor (X10 and X32 and X71) xor (X11 and X30 and X70) xor (X11 and X30 and X72) xor (X11 and X31 and X70) xor (X11 and X32 and X70) xor (X11 and X32 and X71) xor (X12 and X30 and X70) xor (X12 and X30 and X71) xor (X12 and X31 and X70) xor (X12 and X31 and X71) xor (X12 and X32 and X70) xor (X12 and X32 and X72) xor (X20 and X30 and X70) xor (X20 and X30 and X72) xor (X20 and X31 and X71) xor (X20 and X31 and X72) xor (X20 and X32 and X71) xor (X21 and X30 and X70) xor (X21 and X30 and X72) xor (X21 and X31 and X70) xor (X21 and X32 and X70) xor (X21 and X32 and X71) xor (X22 and X30 and X70) xor (X22 and X30 and X71) xor (X22 and X31 and X70) xor (X22 and X31 and X71) xor (X22 and X32 and X70) xor (X22 and X32 and X72) xor (X20 and X40 and X70) xor (X20 and X40 and X72) xor (X20 and X41 and X71) xor (X20 and X41 and X72) xor (X20 and X42 and X71) xor (X21 and X40 and X70) xor (X21 and X40 and X72) xor (X21 and X41 and X70) xor (X21 and X42 and X70) xor (X21 and X42 and X71) xor (X22 and X40 and X70) xor (X22 and X40 and X71) xor (X22 and X41 and X70) xor (X22 and X41 and X71) xor (X22 and X42 and X70) xor (X22 and X42 and X72) xor (X20 and X50 and X70) xor (X20 and X50 and X72) xor (X20 and X51 and X71) xor (X20 and X51 and X72) xor (X20 and X52 and X71) xor (X21 and X50 and X70) xor (X21 and X50 and X72) xor (X21 and X51 and X70) xor (X21 and X52 and X70) xor (X21 and X52 and X71) xor (X22 and X50 and X70) xor (X22 and X50 and X71) xor (X22 and X51 and X70) xor (X22 and X51 and X71) xor (X22 and X52 and X70) xor (X22 and X52 and X72) xor (X10 and X60 and X70) xor (X10 and X60 and X72) xor (X10 and X61 and X71) xor (X10 and X61 and X72) xor (X10 and X62 and X71) xor (X11 and X60 and X70) xor (X11 and X60 and X72) xor (X11 and X61 and X70) xor (X11 and X62 and X70) xor (X11 and X62 and X71) xor (X12 and X60 and X70) xor (X12 and X60 and X71) xor (X12 and X61 and X70) xor (X12 and X61 and X71) xor (X12 and X62 and X70) xor (X12 and X62 and X72) xor (X20 and X60 and X70) xor (X20 and X60 and X72) xor (X20 and X61 and X71) xor (X20 and X61 and X72) xor (X20 and X62 and X71) xor (X21 and X60 and X70) xor (X21 and X60 and X72) xor (X21 and X61 and X70) xor (X21 and X62 and X70) xor (X21 and X62 and X71) xor (X22 and X60 and X70) xor (X22 and X60 and X71) xor (X22 and X61 and X70) xor (X22 and X61 and X71) xor (X22 and X62 and X70) xor (X22 and X62 and X72) xor (X40 and X60 and X70) xor (X40 and X60 and X72) xor (X40 and X61 and X71) xor (X40 and X61 and X72) xor (X40 and X62 and X71) xor (X41 and X60 and X70) xor (X41 and X60 and X72) xor (X41 and X61 and X70) xor (X41 and X62 and X70) xor (X41 and X62 and X71) xor (X42 and X60 and X70) xor (X42 and X60 and X71) xor (X42 and X61 and X70) xor (X42 and X61 and X71) xor (X42 and X62 and X70) xor (X42 and X62 and X72) xor (X50 and X60 and X70) xor (X50 and X60 and X72) xor (X50 and X61 and X71) xor (X50 and X61 and X72) xor (X50 and X62 and X71) xor (X51 and X60 and X70) xor (X51 and X60 and X72) xor (X51 and X61 and X70) xor (X51 and X62 and X70) xor (X51 and X62 and X71) xor (X52 and X60 and X70) xor (X52 and X60 and X71) xor (X52 and X61 and X70) xor (X52 and X61 and X71) xor (X52 and X62 and X70) xor (X52 and X62 and X72));
    F11  <= ((X11) xor (X0_1 and X11) xor (X0_1 and X12) xor (X02 and X11) xor (X0_1 and X13) xor (X0_1 and X21) xor (X0_1 and X22) xor (X02 and X21) xor (X0_1 and X23) xor (X0_1 and X11 and X21) xor (X0_1 and X11 and X22) xor (X0_1 and X12 and X22) xor (X0_1 and X12 and X23) xor (X0_1 and X13 and X22) xor (X02 and X11 and X22) xor (X02 and X11 and X23) xor (X02 and X12 and X21) xor (X02 and X12 and X23) xor (X02 and X13 and X21) xor (X02 and X13 and X22) xor (X03 and X11 and X22) xor (X03 and X12 and X21) xor (X03 and X12 and X23) xor (X03 and X13 and X21) xor (X03 and X13 and X23) xor (X0_1 and X31) xor (X0_1 and X32) xor (X02 and X31) xor (X0_1 and X33) xor (X0_1 and X11 and X31) xor (X0_1 and X11 and X32) xor (X0_1 and X12 and X32) xor (X0_1 and X12 and X33) xor (X0_1 and X13 and X32) xor (X02 and X11 and X32) xor (X02 and X11 and X33) xor (X02 and X12 and X31) xor (X02 and X12 and X33) xor (X02 and X13 and X31) xor (X02 and X13 and X32) xor (X03 and X11 and X32) xor (X03 and X12 and X31) xor (X03 and X12 and X33) xor (X03 and X13 and X31) xor (X03 and X13 and X33) xor (X0_1 and X11 and X41) xor (X0_1 and X11 and X42) xor (X0_1 and X12 and X42) xor (X0_1 and X12 and X43) xor (X0_1 and X13 and X42) xor (X02 and X11 and X42) xor (X02 and X11 and X43) xor (X02 and X12 and X41) xor (X02 and X12 and X43) xor (X02 and X13 and X41) xor (X02 and X13 and X42) xor (X03 and X11 and X42) xor (X03 and X12 and X41) xor (X03 and X12 and X43) xor (X03 and X13 and X41) xor (X03 and X13 and X43) xor (X21 and X41) xor (X21 and X42) xor (X22 and X41) xor (X21 and X43) xor (X0_1 and X21 and X41) xor (X0_1 and X21 and X42) xor (X0_1 and X22 and X42) xor (X0_1 and X22 and X43) xor (X0_1 and X23 and X42) xor (X02 and X21 and X42) xor (X02 and X21 and X43) xor (X02 and X22 and X41) xor (X02 and X22 and X43) xor (X02 and X23 and X41) xor (X02 and X23 and X42) xor (X03 and X21 and X42) xor (X03 and X22 and X41) xor (X03 and X22 and X43) xor (X03 and X23 and X41) xor (X03 and X23 and X43) xor (X0_1 and X31 and X41) xor (X0_1 and X31 and X42) xor (X0_1 and X32 and X42) xor (X0_1 and X32 and X43) xor (X0_1 and X33 and X42) xor (X02 and X31 and X42) xor (X02 and X31 and X43) xor (X02 and X32 and X41) xor (X02 and X32 and X43) xor (X02 and X33 and X41) xor (X02 and X33 and X42) xor (X03 and X31 and X42) xor (X03 and X32 and X41) xor (X03 and X32 and X43) xor (X03 and X33 and X41) xor (X03 and X33 and X43) xor (X51) xor (X11 and X51) xor (X11 and X52) xor (X12 and X51) xor (X11 and X53) xor (X21 and X51) xor (X21 and X52) xor (X22 and X51) xor (X21 and X53) xor (X31 and X51) xor (X31 and X52) xor (X32 and X51) xor (X31 and X53) xor (X11 and X31 and X51) xor (X11 and X31 and X52) xor (X11 and X32 and X52) xor (X11 and X32 and X53) xor (X11 and X33 and X52) xor (X12 and X31 and X52) xor (X12 and X31 and X53) xor (X12 and X32 and X51) xor (X12 and X32 and X53) xor (X12 and X33 and X51) xor (X12 and X33 and X52) xor (X13 and X31 and X52) xor (X13 and X32 and X51) xor (X13 and X32 and X53) xor (X13 and X33 and X51) xor (X13 and X33 and X53) xor (X21 and X31 and X51) xor (X21 and X31 and X52) xor (X21 and X32 and X52) xor (X21 and X32 and X53) xor (X21 and X33 and X52) xor (X22 and X31 and X52) xor (X22 and X31 and X53) xor (X22 and X32 and X51) xor (X22 and X32 and X53) xor (X22 and X33 and X51) xor (X22 and X33 and X52) xor (X23 and X31 and X52) xor (X23 and X32 and X51) xor (X23 and X32 and X53) xor (X23 and X33 and X51) xor (X23 and X33 and X53) xor (X31 and X41 and X51) xor (X31 and X41 and X52) xor (X31 and X42 and X52) xor (X31 and X42 and X53) xor (X31 and X43 and X52) xor (X32 and X41 and X52) xor (X32 and X41 and X53) xor (X32 and X42 and X51) xor (X32 and X42 and X53) xor (X32 and X43 and X51) xor (X32 and X43 and X52) xor (X33 and X41 and X52) xor (X33 and X42 and X51) xor (X33 and X42 and X53) xor (X33 and X43 and X51) xor (X33 and X43 and X53) xor (X61) xor (X11 and X61) xor (X11 and X62) xor (X12 and X61) xor (X11 and X63) xor (X0_1 and X11 and X61) xor (X0_1 and X11 and X62) xor (X0_1 and X12 and X62) xor (X0_1 and X12 and X63) xor (X0_1 and X13 and X62) xor (X02 and X11 and X62) xor (X02 and X11 and X63) xor (X02 and X12 and X61) xor (X02 and X12 and X63) xor (X02 and X13 and X61) xor (X02 and X13 and X62) xor (X03 and X11 and X62) xor (X03 and X12 and X61) xor (X03 and X12 and X63) xor (X03 and X13 and X61) xor (X03 and X13 and X63) xor (X21 and X61) xor (X21 and X62) xor (X22 and X61) xor (X21 and X63) xor (X0_1 and X21 and X61) xor (X0_1 and X21 and X62) xor (X0_1 and X22 and X62) xor (X0_1 and X22 and X63) xor (X0_1 and X23 and X62) xor (X02 and X21 and X62) xor (X02 and X21 and X63) xor (X02 and X22 and X61) xor (X02 and X22 and X63) xor (X02 and X23 and X61) xor (X02 and X23 and X62) xor (X03 and X21 and X62) xor (X03 and X22 and X61) xor (X03 and X22 and X63) xor (X03 and X23 and X61) xor (X03 and X23 and X63) xor (X0_1 and X31 and X61) xor (X0_1 and X31 and X62) xor (X0_1 and X32 and X62) xor (X0_1 and X32 and X63) xor (X0_1 and X33 and X62) xor (X02 and X31 and X62) xor (X02 and X31 and X63) xor (X02 and X32 and X61) xor (X02 and X32 and X63) xor (X02 and X33 and X61) xor (X02 and X33 and X62) xor (X03 and X31 and X62) xor (X03 and X32 and X61) xor (X03 and X32 and X63) xor (X03 and X33 and X61) xor (X03 and X33 and X63) xor (X41 and X61) xor (X41 and X62) xor (X42 and X61) xor (X41 and X63) xor (X11 and X41 and X61) xor (X11 and X41 and X62) xor (X11 and X42 and X62) xor (X11 and X42 and X63) xor (X11 and X43 and X62) xor (X12 and X41 and X62) xor (X12 and X41 and X63) xor (X12 and X42 and X61) xor (X12 and X42 and X63) xor (X12 and X43 and X61) xor (X12 and X43 and X62) xor (X13 and X41 and X62) xor (X13 and X42 and X61) xor (X13 and X42 and X63) xor (X13 and X43 and X61) xor (X13 and X43 and X63) xor (X31 and X51 and X61) xor (X31 and X51 and X62) xor (X31 and X52 and X62) xor (X31 and X52 and X63) xor (X31 and X53 and X62) xor (X32 and X51 and X62) xor (X32 and X51 and X63) xor (X32 and X52 and X61) xor (X32 and X52 and X63) xor (X32 and X53 and X61) xor (X32 and X53 and X62) xor (X33 and X51 and X62) xor (X33 and X52 and X61) xor (X33 and X52 and X63) xor (X33 and X53 and X61) xor (X33 and X53 and X63) xor (X41 and X51 and X61) xor (X41 and X51 and X62) xor (X41 and X52 and X62) xor (X41 and X52 and X63) xor (X41 and X53 and X62) xor (X42 and X51 and X62) xor (X42 and X51 and X63) xor (X42 and X52 and X61) xor (X42 and X52 and X63) xor (X42 and X53 and X61) xor (X42 and X53 and X62) xor (X43 and X51 and X62) xor (X43 and X52 and X61) xor (X43 and X52 and X63) xor (X43 and X53 and X61) xor (X43 and X53 and X63) xor (X71) xor (X11 and X71) xor (X11 and X72) xor (X12 and X71) xor (X11 and X73) xor (X0_1 and X11 and X71) xor (X0_1 and X11 and X72) xor (X0_1 and X12 and X72) xor (X0_1 and X12 and X73) xor (X0_1 and X13 and X72) xor (X02 and X11 and X72) xor (X02 and X11 and X73) xor (X02 and X12 and X71) xor (X02 and X12 and X73) xor (X02 and X13 and X71) xor (X02 and X13 and X72) xor (X03 and X11 and X72) xor (X03 and X12 and X71) xor (X03 and X12 and X73) xor (X03 and X13 and X71) xor (X03 and X13 and X73) xor (X0_1 and X21 and X71) xor (X0_1 and X21 and X72) xor (X0_1 and X22 and X72) xor (X0_1 and X22 and X73) xor (X0_1 and X23 and X72) xor (X02 and X21 and X72) xor (X02 and X21 and X73) xor (X02 and X22 and X71) xor (X02 and X22 and X73) xor (X02 and X23 and X71) xor (X02 and X23 and X72) xor (X03 and X21 and X72) xor (X03 and X22 and X71) xor (X03 and X22 and X73) xor (X03 and X23 and X71) xor (X03 and X23 and X73) xor (X0_1 and X31 and X71) xor (X0_1 and X31 and X72) xor (X0_1 and X32 and X72) xor (X0_1 and X32 and X73) xor (X0_1 and X33 and X72) xor (X02 and X31 and X72) xor (X02 and X31 and X73) xor (X02 and X32 and X71) xor (X02 and X32 and X73) xor (X02 and X33 and X71) xor (X02 and X33 and X72) xor (X03 and X31 and X72) xor (X03 and X32 and X71) xor (X03 and X32 and X73) xor (X03 and X33 and X71) xor (X03 and X33 and X73) xor (X11 and X31 and X71) xor (X11 and X31 and X72) xor (X11 and X32 and X72) xor (X11 and X32 and X73) xor (X11 and X33 and X72) xor (X12 and X31 and X72) xor (X12 and X31 and X73) xor (X12 and X32 and X71) xor (X12 and X32 and X73) xor (X12 and X33 and X71) xor (X12 and X33 and X72) xor (X13 and X31 and X72) xor (X13 and X32 and X71) xor (X13 and X32 and X73) xor (X13 and X33 and X71) xor (X13 and X33 and X73) xor (X21 and X31 and X71) xor (X21 and X31 and X72) xor (X21 and X32 and X72) xor (X21 and X32 and X73) xor (X21 and X33 and X72) xor (X22 and X31 and X72) xor (X22 and X31 and X73) xor (X22 and X32 and X71) xor (X22 and X32 and X73) xor (X22 and X33 and X71) xor (X22 and X33 and X72) xor (X23 and X31 and X72) xor (X23 and X32 and X71) xor (X23 and X32 and X73) xor (X23 and X33 and X71) xor (X23 and X33 and X73) xor (X21 and X41 and X71) xor (X21 and X41 and X72) xor (X21 and X42 and X72) xor (X21 and X42 and X73) xor (X21 and X43 and X72) xor (X22 and X41 and X72) xor (X22 and X41 and X73) xor (X22 and X42 and X71) xor (X22 and X42 and X73) xor (X22 and X43 and X71) xor (X22 and X43 and X72) xor (X23 and X41 and X72) xor (X23 and X42 and X71) xor (X23 and X42 and X73) xor (X23 and X43 and X71) xor (X23 and X43 and X73) xor (X21 and X51 and X71) xor (X21 and X51 and X72) xor (X21 and X52 and X72) xor (X21 and X52 and X73) xor (X21 and X53 and X72) xor (X22 and X51 and X72) xor (X22 and X51 and X73) xor (X22 and X52 and X71) xor (X22 and X52 and X73) xor (X22 and X53 and X71) xor (X22 and X53 and X72) xor (X23 and X51 and X72) xor (X23 and X52 and X71) xor (X23 and X52 and X73) xor (X23 and X53 and X71) xor (X23 and X53 and X73) xor (X11 and X61 and X71) xor (X11 and X61 and X72) xor (X11 and X62 and X72) xor (X11 and X62 and X73) xor (X11 and X63 and X72) xor (X12 and X61 and X72) xor (X12 and X61 and X73) xor (X12 and X62 and X71) xor (X12 and X62 and X73) xor (X12 and X63 and X71) xor (X12 and X63 and X72) xor (X13 and X61 and X72) xor (X13 and X62 and X71) xor (X13 and X62 and X73) xor (X13 and X63 and X71) xor (X13 and X63 and X73) xor (X21 and X61 and X71) xor (X21 and X61 and X72) xor (X21 and X62 and X72) xor (X21 and X62 and X73) xor (X21 and X63 and X72) xor (X22 and X61 and X72) xor (X22 and X61 and X73) xor (X22 and X62 and X71) xor (X22 and X62 and X73) xor (X22 and X63 and X71) xor (X22 and X63 and X72) xor (X23 and X61 and X72) xor (X23 and X62 and X71) xor (X23 and X62 and X73) xor (X23 and X63 and X71) xor (X23 and X63 and X73) xor (X41 and X61 and X71) xor (X41 and X61 and X72) xor (X41 and X62 and X72) xor (X41 and X62 and X73) xor (X41 and X63 and X72) xor (X42 and X61 and X72) xor (X42 and X61 and X73) xor (X42 and X62 and X71) xor (X42 and X62 and X73) xor (X42 and X63 and X71) xor (X42 and X63 and X72) xor (X43 and X61 and X72) xor (X43 and X62 and X71) xor (X43 and X62 and X73) xor (X43 and X63 and X71) xor (X43 and X63 and X73) xor (X51 and X61 and X71) xor (X51 and X61 and X72) xor (X51 and X62 and X72) xor (X51 and X62 and X73) xor (X51 and X63 and X72) xor (X52 and X61 and X72) xor (X52 and X61 and X73) xor (X52 and X62 and X71) xor (X52 and X62 and X73) xor (X52 and X63 and X71) xor (X52 and X63 and X72) xor (X53 and X61 and X72) xor (X53 and X62 and X71) xor (X53 and X62 and X73) xor (X53 and X63 and X71) xor (X53 and X63 and X73));
    F12  <= ((X12) xor (X02 and X12) xor (X00 and X13) xor (X02 and X13) xor (X03 and X12) xor (X02 and X22) xor (X00 and X23) xor (X02 and X23) xor (X03 and X22) xor (X00 and X10 and X23) xor (X00 and X12 and X20) xor (X00 and X12 and X22) xor (X00 and X12 and X23) xor (X00 and X13 and X20) xor (X00 and X13 and X22) xor (X02 and X10 and X22) xor (X02 and X10 and X23) xor (X02 and X13 and X20) xor (X02 and X13 and X23) xor (X03 and X10 and X20) xor (X03 and X10 and X22) xor (X03 and X10 and X23) xor (X03 and X12 and X20) xor (X03 and X12 and X22) xor (X03 and X13 and X22) xor (X02 and X32) xor (X00 and X33) xor (X02 and X33) xor (X03 and X32) xor (X00 and X10 and X33) xor (X00 and X12 and X30) xor (X00 and X12 and X32) xor (X00 and X12 and X33) xor (X00 and X13 and X30) xor (X00 and X13 and X32) xor (X02 and X10 and X32) xor (X02 and X10 and X33) xor (X02 and X13 and X30) xor (X02 and X13 and X33) xor (X03 and X10 and X30) xor (X03 and X10 and X32) xor (X03 and X10 and X33) xor (X03 and X12 and X30) xor (X03 and X12 and X32) xor (X03 and X13 and X32) xor (X00 and X10 and X43) xor (X00 and X12 and X40) xor (X00 and X12 and X42) xor (X00 and X12 and X43) xor (X00 and X13 and X40) xor (X00 and X13 and X42) xor (X02 and X10 and X42) xor (X02 and X10 and X43) xor (X02 and X13 and X40) xor (X02 and X13 and X43) xor (X03 and X10 and X40) xor (X03 and X10 and X42) xor (X03 and X10 and X43) xor (X03 and X12 and X40) xor (X03 and X12 and X42) xor (X03 and X13 and X42) xor (X22 and X42) xor (X20 and X43) xor (X22 and X43) xor (X23 and X42) xor (X00 and X20 and X43) xor (X00 and X22 and X40) xor (X00 and X22 and X42) xor (X00 and X22 and X43) xor (X00 and X23 and X40) xor (X00 and X23 and X42) xor (X02 and X20 and X42) xor (X02 and X20 and X43) xor (X02 and X23 and X40) xor (X02 and X23 and X43) xor (X03 and X20 and X40) xor (X03 and X20 and X42) xor (X03 and X20 and X43) xor (X03 and X22 and X40) xor (X03 and X22 and X42) xor (X03 and X23 and X42) xor (X00 and X30 and X43) xor (X00 and X32 and X40) xor (X00 and X32 and X42) xor (X00 and X32 and X43) xor (X00 and X33 and X40) xor (X00 and X33 and X42) xor (X02 and X30 and X42) xor (X02 and X30 and X43) xor (X02 and X33 and X40) xor (X02 and X33 and X43) xor (X03 and X30 and X40) xor (X03 and X30 and X42) xor (X03 and X30 and X43) xor (X03 and X32 and X40) xor (X03 and X32 and X42) xor (X03 and X33 and X42) xor (X52) xor (X12 and X52) xor (X10 and X53) xor (X12 and X53) xor (X13 and X52) xor (X22 and X52) xor (X20 and X53) xor (X22 and X53) xor (X23 and X52) xor (X32 and X52) xor (X30 and X53) xor (X32 and X53) xor (X33 and X52) xor (X10 and X30 and X53) xor (X10 and X32 and X50) xor (X10 and X32 and X52) xor (X10 and X32 and X53) xor (X10 and X33 and X50) xor (X10 and X33 and X52) xor (X12 and X30 and X52) xor (X12 and X30 and X53) xor (X12 and X33 and X50) xor (X12 and X33 and X53) xor (X13 and X30 and X50) xor (X13 and X30 and X52) xor (X13 and X30 and X53) xor (X13 and X32 and X50) xor (X13 and X32 and X52) xor (X13 and X33 and X52) xor (X20 and X30 and X53) xor (X20 and X32 and X50) xor (X20 and X32 and X52) xor (X20 and X32 and X53) xor (X20 and X33 and X50) xor (X20 and X33 and X52) xor (X22 and X30 and X52) xor (X22 and X30 and X53) xor (X22 and X33 and X50) xor (X22 and X33 and X53) xor (X23 and X30 and X50) xor (X23 and X30 and X52) xor (X23 and X30 and X53) xor (X23 and X32 and X50) xor (X23 and X32 and X52) xor (X23 and X33 and X52) xor (X30 and X40 and X53) xor (X30 and X42 and X50) xor (X30 and X42 and X52) xor (X30 and X42 and X53) xor (X30 and X43 and X50) xor (X30 and X43 and X52) xor (X32 and X40 and X52) xor (X32 and X40 and X53) xor (X32 and X43 and X50) xor (X32 and X43 and X53) xor (X33 and X40 and X50) xor (X33 and X40 and X52) xor (X33 and X40 and X53) xor (X33 and X42 and X50) xor (X33 and X42 and X52) xor (X33 and X43 and X52) xor (X62) xor (X12 and X62) xor (X10 and X63) xor (X12 and X63) xor (X13 and X62) xor (X00 and X10 and X63) xor (X00 and X12 and X60) xor (X00 and X12 and X62) xor (X00 and X12 and X63) xor (X00 and X13 and X60) xor (X00 and X13 and X62) xor (X02 and X10 and X62) xor (X02 and X10 and X63) xor (X02 and X13 and X60) xor (X02 and X13 and X63) xor (X03 and X10 and X60) xor (X03 and X10 and X62) xor (X03 and X10 and X63) xor (X03 and X12 and X60) xor (X03 and X12 and X62) xor (X03 and X13 and X62) xor (X22 and X62) xor (X20 and X63) xor (X22 and X63) xor (X23 and X62) xor (X00 and X20 and X63) xor (X00 and X22 and X60) xor (X00 and X22 and X62) xor (X00 and X22 and X63) xor (X00 and X23 and X60) xor (X00 and X23 and X62) xor (X02 and X20 and X62) xor (X02 and X20 and X63) xor (X02 and X23 and X60) xor (X02 and X23 and X63) xor (X03 and X20 and X60) xor (X03 and X20 and X62) xor (X03 and X20 and X63) xor (X03 and X22 and X60) xor (X03 and X22 and X62) xor (X03 and X23 and X62) xor (X00 and X30 and X63) xor (X00 and X32 and X60) xor (X00 and X32 and X62) xor (X00 and X32 and X63) xor (X00 and X33 and X60) xor (X00 and X33 and X62) xor (X02 and X30 and X62) xor (X02 and X30 and X63) xor (X02 and X33 and X60) xor (X02 and X33 and X63) xor (X03 and X30 and X60) xor (X03 and X30 and X62) xor (X03 and X30 and X63) xor (X03 and X32 and X60) xor (X03 and X32 and X62) xor (X03 and X33 and X62) xor (X42 and X62) xor (X40 and X63) xor (X42 and X63) xor (X43 and X62) xor (X10 and X40 and X63) xor (X10 and X42 and X60) xor (X10 and X42 and X62) xor (X10 and X42 and X63) xor (X10 and X43 and X60) xor (X10 and X43 and X62) xor (X12 and X40 and X62) xor (X12 and X40 and X63) xor (X12 and X43 and X60) xor (X12 and X43 and X63) xor (X13 and X40 and X60) xor (X13 and X40 and X62) xor (X13 and X40 and X63) xor (X13 and X42 and X60) xor (X13 and X42 and X62) xor (X13 and X43 and X62) xor (X30 and X50 and X63) xor (X30 and X52 and X60) xor (X30 and X52 and X62) xor (X30 and X52 and X63) xor (X30 and X53 and X60) xor (X30 and X53 and X62) xor (X32 and X50 and X62) xor (X32 and X50 and X63) xor (X32 and X53 and X60) xor (X32 and X53 and X63) xor (X33 and X50 and X60) xor (X33 and X50 and X62) xor (X33 and X50 and X63) xor (X33 and X52 and X60) xor (X33 and X52 and X62) xor (X33 and X53 and X62) xor (X40 and X50 and X63) xor (X40 and X52 and X60) xor (X40 and X52 and X62) xor (X40 and X52 and X63) xor (X40 and X53 and X60) xor (X40 and X53 and X62) xor (X42 and X50 and X62) xor (X42 and X50 and X63) xor (X42 and X53 and X60) xor (X42 and X53 and X63) xor (X43 and X50 and X60) xor (X43 and X50 and X62) xor (X43 and X50 and X63) xor (X43 and X52 and X60) xor (X43 and X52 and X62) xor (X43 and X53 and X62) xor (X72) xor (X12 and X72) xor (X10 and X73) xor (X12 and X73) xor (X13 and X72) xor (X00 and X10 and X73) xor (X00 and X12 and X70) xor (X00 and X12 and X72) xor (X00 and X12 and X73) xor (X00 and X13 and X70) xor (X00 and X13 and X72) xor (X02 and X10 and X72) xor (X02 and X10 and X73) xor (X02 and X13 and X70) xor (X02 and X13 and X73) xor (X03 and X10 and X70) xor (X03 and X10 and X72) xor (X03 and X10 and X73) xor (X03 and X12 and X70) xor (X03 and X12 and X72) xor (X03 and X13 and X72) xor (X00 and X20 and X73) xor (X00 and X22 and X70) xor (X00 and X22 and X72) xor (X00 and X22 and X73) xor (X00 and X23 and X70) xor (X00 and X23 and X72) xor (X02 and X20 and X72) xor (X02 and X20 and X73) xor (X02 and X23 and X70) xor (X02 and X23 and X73) xor (X03 and X20 and X70) xor (X03 and X20 and X72) xor (X03 and X20 and X73) xor (X03 and X22 and X70) xor (X03 and X22 and X72) xor (X03 and X23 and X72) xor (X00 and X30 and X73) xor (X00 and X32 and X70) xor (X00 and X32 and X72) xor (X00 and X32 and X73) xor (X00 and X33 and X70) xor (X00 and X33 and X72) xor (X02 and X30 and X72) xor (X02 and X30 and X73) xor (X02 and X33 and X70) xor (X02 and X33 and X73) xor (X03 and X30 and X70) xor (X03 and X30 and X72) xor (X03 and X30 and X73) xor (X03 and X32 and X70) xor (X03 and X32 and X72) xor (X03 and X33 and X72) xor (X10 and X30 and X73) xor (X10 and X32 and X70) xor (X10 and X32 and X72) xor (X10 and X32 and X73) xor (X10 and X33 and X70) xor (X10 and X33 and X72) xor (X12 and X30 and X72) xor (X12 and X30 and X73) xor (X12 and X33 and X70) xor (X12 and X33 and X73) xor (X13 and X30 and X70) xor (X13 and X30 and X72) xor (X13 and X30 and X73) xor (X13 and X32 and X70) xor (X13 and X32 and X72) xor (X13 and X33 and X72) xor (X20 and X30 and X73) xor (X20 and X32 and X70) xor (X20 and X32 and X72) xor (X20 and X32 and X73) xor (X20 and X33 and X70) xor (X20 and X33 and X72) xor (X22 and X30 and X72) xor (X22 and X30 and X73) xor (X22 and X33 and X70) xor (X22 and X33 and X73) xor (X23 and X30 and X70) xor (X23 and X30 and X72) xor (X23 and X30 and X73) xor (X23 and X32 and X70) xor (X23 and X32 and X72) xor (X23 and X33 and X72) xor (X20 and X40 and X73) xor (X20 and X42 and X70) xor (X20 and X42 and X72) xor (X20 and X42 and X73) xor (X20 and X43 and X70) xor (X20 and X43 and X72) xor (X22 and X40 and X72) xor (X22 and X40 and X73) xor (X22 and X43 and X70) xor (X22 and X43 and X73) xor (X23 and X40 and X70) xor (X23 and X40 and X72) xor (X23 and X40 and X73) xor (X23 and X42 and X70) xor (X23 and X42 and X72) xor (X23 and X43 and X72) xor (X20 and X50 and X73) xor (X20 and X52 and X70) xor (X20 and X52 and X72) xor (X20 and X52 and X73) xor (X20 and X53 and X70) xor (X20 and X53 and X72) xor (X22 and X50 and X72) xor (X22 and X50 and X73) xor (X22 and X53 and X70) xor (X22 and X53 and X73) xor (X23 and X50 and X70) xor (X23 and X50 and X72) xor (X23 and X50 and X73) xor (X23 and X52 and X70) xor (X23 and X52 and X72) xor (X23 and X53 and X72) xor (X10 and X60 and X73) xor (X10 and X62 and X70) xor (X10 and X62 and X72) xor (X10 and X62 and X73) xor (X10 and X63 and X70) xor (X10 and X63 and X72) xor (X12 and X60 and X72) xor (X12 and X60 and X73) xor (X12 and X63 and X70) xor (X12 and X63 and X73) xor (X13 and X60 and X70) xor (X13 and X60 and X72) xor (X13 and X60 and X73) xor (X13 and X62 and X70) xor (X13 and X62 and X72) xor (X13 and X63 and X72) xor (X20 and X60 and X73) xor (X20 and X62 and X70) xor (X20 and X62 and X72) xor (X20 and X62 and X73) xor (X20 and X63 and X70) xor (X20 and X63 and X72) xor (X22 and X60 and X72) xor (X22 and X60 and X73) xor (X22 and X63 and X70) xor (X22 and X63 and X73) xor (X23 and X60 and X70) xor (X23 and X60 and X72) xor (X23 and X60 and X73) xor (X23 and X62 and X70) xor (X23 and X62 and X72) xor (X23 and X63 and X72) xor (X40 and X60 and X73) xor (X40 and X62 and X70) xor (X40 and X62 and X72) xor (X40 and X62 and X73) xor (X40 and X63 and X70) xor (X40 and X63 and X72) xor (X42 and X60 and X72) xor (X42 and X60 and X73) xor (X42 and X63 and X70) xor (X42 and X63 and X73) xor (X43 and X60 and X70) xor (X43 and X60 and X72) xor (X43 and X60 and X73) xor (X43 and X62 and X70) xor (X43 and X62 and X72) xor (X43 and X63 and X72) xor (X50 and X60 and X73) xor (X50 and X62 and X70) xor (X50 and X62 and X72) xor (X50 and X62 and X73) xor (X50 and X63 and X70) xor (X50 and X63 and X72) xor (X52 and X60 and X72) xor (X52 and X60 and X73) xor (X52 and X63 and X70) xor (X52 and X63 and X73) xor (X53 and X60 and X70) xor (X53 and X60 and X72) xor (X53 and X60 and X73) xor (X53 and X62 and X70) xor (X53 and X62 and X72) xor (X53 and X63 and X72));
    F13  <= ((X13) xor (X03 and X13) xor (X03 and X10) xor (X03 and X11) xor (X0_1 and X10) xor (X03 and X23) xor (X03 and X20) xor (X03 and X21) xor (X0_1 and X20) xor (X00 and X10 and X21) xor (X00 and X11 and X20) xor (X00 and X11 and X23) xor (X00 and X13 and X21) xor (X00 and X13 and X23) xor (X0_1 and X10 and X21) xor (X0_1 and X10 and X23) xor (X0_1 and X11 and X23) xor (X0_1 and X13 and X20) xor (X0_1 and X13 and X21) xor (X0_1 and X13 and X23) xor (X03 and X10 and X21) xor (X03 and X11 and X20) xor (X03 and X11 and X21) xor (X03 and X11 and X23) xor (X03 and X13 and X20) xor (X03 and X33) xor (X03 and X30) xor (X03 and X31) xor (X0_1 and X30) xor (X00 and X10 and X31) xor (X00 and X11 and X30) xor (X00 and X11 and X33) xor (X00 and X13 and X31) xor (X00 and X13 and X33) xor (X0_1 and X10 and X31) xor (X0_1 and X10 and X33) xor (X0_1 and X11 and X33) xor (X0_1 and X13 and X30) xor (X0_1 and X13 and X31) xor (X0_1 and X13 and X33) xor (X03 and X10 and X31) xor (X03 and X11 and X30) xor (X03 and X11 and X31) xor (X03 and X11 and X33) xor (X03 and X13 and X30) xor (X00 and X10 and X41) xor (X00 and X11 and X40) xor (X00 and X11 and X43) xor (X00 and X13 and X41) xor (X00 and X13 and X43) xor (X0_1 and X10 and X41) xor (X0_1 and X10 and X43) xor (X0_1 and X11 and X43) xor (X0_1 and X13 and X40) xor (X0_1 and X13 and X41) xor (X0_1 and X13 and X43) xor (X03 and X10 and X41) xor (X03 and X11 and X40) xor (X03 and X11 and X41) xor (X03 and X11 and X43) xor (X03 and X13 and X40) xor (X23 and X43) xor (X23 and X40) xor (X23 and X41) xor (X21 and X40) xor (X00 and X20 and X41) xor (X00 and X21 and X40) xor (X00 and X21 and X43) xor (X00 and X23 and X41) xor (X00 and X23 and X43) xor (X0_1 and X20 and X41) xor (X0_1 and X20 and X43) xor (X0_1 and X21 and X43) xor (X0_1 and X23 and X40) xor (X0_1 and X23 and X41) xor (X0_1 and X23 and X43) xor (X03 and X20 and X41) xor (X03 and X21 and X40) xor (X03 and X21 and X41) xor (X03 and X21 and X43) xor (X03 and X23 and X40) xor (X00 and X30 and X41) xor (X00 and X31 and X40) xor (X00 and X31 and X43) xor (X00 and X33 and X41) xor (X00 and X33 and X43) xor (X0_1 and X30 and X41) xor (X0_1 and X30 and X43) xor (X0_1 and X31 and X43) xor (X0_1 and X33 and X40) xor (X0_1 and X33 and X41) xor (X0_1 and X33 and X43) xor (X03 and X30 and X41) xor (X03 and X31 and X40) xor (X03 and X31 and X41) xor (X03 and X31 and X43) xor (X03 and X33 and X40) xor (X53) xor (X13 and X53) xor (X13 and X50) xor (X13 and X51) xor (X11 and X50) xor (X23 and X53) xor (X23 and X50) xor (X23 and X51) xor (X21 and X50) xor (X33 and X53) xor (X33 and X50) xor (X33 and X51) xor (X31 and X50) xor (X10 and X30 and X51) xor (X10 and X31 and X50) xor (X10 and X31 and X53) xor (X10 and X33 and X51) xor (X10 and X33 and X53) xor (X11 and X30 and X51) xor (X11 and X30 and X53) xor (X11 and X31 and X53) xor (X11 and X33 and X50) xor (X11 and X33 and X51) xor (X11 and X33 and X53) xor (X13 and X30 and X51) xor (X13 and X31 and X50) xor (X13 and X31 and X51) xor (X13 and X31 and X53) xor (X13 and X33 and X50) xor (X20 and X30 and X51) xor (X20 and X31 and X50) xor (X20 and X31 and X53) xor (X20 and X33 and X51) xor (X20 and X33 and X53) xor (X21 and X30 and X51) xor (X21 and X30 and X53) xor (X21 and X31 and X53) xor (X21 and X33 and X50) xor (X21 and X33 and X51) xor (X21 and X33 and X53) xor (X23 and X30 and X51) xor (X23 and X31 and X50) xor (X23 and X31 and X51) xor (X23 and X31 and X53) xor (X23 and X33 and X50) xor (X30 and X40 and X51) xor (X30 and X41 and X50) xor (X30 and X41 and X53) xor (X30 and X43 and X51) xor (X30 and X43 and X53) xor (X31 and X40 and X51) xor (X31 and X40 and X53) xor (X31 and X41 and X53) xor (X31 and X43 and X50) xor (X31 and X43 and X51) xor (X31 and X43 and X53) xor (X33 and X40 and X51) xor (X33 and X41 and X50) xor (X33 and X41 and X51) xor (X33 and X41 and X53) xor (X33 and X43 and X50) xor (X63) xor (X13 and X63) xor (X13 and X60) xor (X13 and X61) xor (X11 and X60) xor (X00 and X10 and X61) xor (X00 and X11 and X60) xor (X00 and X11 and X63) xor (X00 and X13 and X61) xor (X00 and X13 and X63) xor (X0_1 and X10 and X61) xor (X0_1 and X10 and X63) xor (X0_1 and X11 and X63) xor (X0_1 and X13 and X60) xor (X0_1 and X13 and X61) xor (X0_1 and X13 and X63) xor (X03 and X10 and X61) xor (X03 and X11 and X60) xor (X03 and X11 and X61) xor (X03 and X11 and X63) xor (X03 and X13 and X60) xor (X23 and X63) xor (X23 and X60) xor (X23 and X61) xor (X21 and X60) xor (X00 and X20 and X61) xor (X00 and X21 and X60) xor (X00 and X21 and X63) xor (X00 and X23 and X61) xor (X00 and X23 and X63) xor (X0_1 and X20 and X61) xor (X0_1 and X20 and X63) xor (X0_1 and X21 and X63) xor (X0_1 and X23 and X60) xor (X0_1 and X23 and X61) xor (X0_1 and X23 and X63) xor (X03 and X20 and X61) xor (X03 and X21 and X60) xor (X03 and X21 and X61) xor (X03 and X21 and X63) xor (X03 and X23 and X60) xor (X00 and X30 and X61) xor (X00 and X31 and X60) xor (X00 and X31 and X63) xor (X00 and X33 and X61) xor (X00 and X33 and X63) xor (X0_1 and X30 and X61) xor (X0_1 and X30 and X63) xor (X0_1 and X31 and X63) xor (X0_1 and X33 and X60) xor (X0_1 and X33 and X61) xor (X0_1 and X33 and X63) xor (X03 and X30 and X61) xor (X03 and X31 and X60) xor (X03 and X31 and X61) xor (X03 and X31 and X63) xor (X03 and X33 and X60) xor (X43 and X63) xor (X43 and X60) xor (X43 and X61) xor (X41 and X60) xor (X10 and X40 and X61) xor (X10 and X41 and X60) xor (X10 and X41 and X63) xor (X10 and X43 and X61) xor (X10 and X43 and X63) xor (X11 and X40 and X61) xor (X11 and X40 and X63) xor (X11 and X41 and X63) xor (X11 and X43 and X60) xor (X11 and X43 and X61) xor (X11 and X43 and X63) xor (X13 and X40 and X61) xor (X13 and X41 and X60) xor (X13 and X41 and X61) xor (X13 and X41 and X63) xor (X13 and X43 and X60) xor (X30 and X50 and X61) xor (X30 and X51 and X60) xor (X30 and X51 and X63) xor (X30 and X53 and X61) xor (X30 and X53 and X63) xor (X31 and X50 and X61) xor (X31 and X50 and X63) xor (X31 and X51 and X63) xor (X31 and X53 and X60) xor (X31 and X53 and X61) xor (X31 and X53 and X63) xor (X33 and X50 and X61) xor (X33 and X51 and X60) xor (X33 and X51 and X61) xor (X33 and X51 and X63) xor (X33 and X53 and X60) xor (X40 and X50 and X61) xor (X40 and X51 and X60) xor (X40 and X51 and X63) xor (X40 and X53 and X61) xor (X40 and X53 and X63) xor (X41 and X50 and X61) xor (X41 and X50 and X63) xor (X41 and X51 and X63) xor (X41 and X53 and X60) xor (X41 and X53 and X61) xor (X41 and X53 and X63) xor (X43 and X50 and X61) xor (X43 and X51 and X60) xor (X43 and X51 and X61) xor (X43 and X51 and X63) xor (X43 and X53 and X60) xor (X73) xor (X13 and X73) xor (X13 and X70) xor (X13 and X71) xor (X11 and X70) xor (X00 and X10 and X71) xor (X00 and X11 and X70) xor (X00 and X11 and X73) xor (X00 and X13 and X71) xor (X00 and X13 and X73) xor (X0_1 and X10 and X71) xor (X0_1 and X10 and X73) xor (X0_1 and X11 and X73) xor (X0_1 and X13 and X70) xor (X0_1 and X13 and X71) xor (X0_1 and X13 and X73) xor (X03 and X10 and X71) xor (X03 and X11 and X70) xor (X03 and X11 and X71) xor (X03 and X11 and X73) xor (X03 and X13 and X70) xor (X00 and X20 and X71) xor (X00 and X21 and X70) xor (X00 and X21 and X73) xor (X00 and X23 and X71) xor (X00 and X23 and X73) xor (X0_1 and X20 and X71) xor (X0_1 and X20 and X73) xor (X0_1 and X21 and X73) xor (X0_1 and X23 and X70) xor (X0_1 and X23 and X71) xor (X0_1 and X23 and X73) xor (X03 and X20 and X71) xor (X03 and X21 and X70) xor (X03 and X21 and X71) xor (X03 and X21 and X73) xor (X03 and X23 and X70) xor (X00 and X30 and X71) xor (X00 and X31 and X70) xor (X00 and X31 and X73) xor (X00 and X33 and X71) xor (X00 and X33 and X73) xor (X0_1 and X30 and X71) xor (X0_1 and X30 and X73) xor (X0_1 and X31 and X73) xor (X0_1 and X33 and X70) xor (X0_1 and X33 and X71) xor (X0_1 and X33 and X73) xor (X03 and X30 and X71) xor (X03 and X31 and X70) xor (X03 and X31 and X71) xor (X03 and X31 and X73) xor (X03 and X33 and X70) xor (X10 and X30 and X71) xor (X10 and X31 and X70) xor (X10 and X31 and X73) xor (X10 and X33 and X71) xor (X10 and X33 and X73) xor (X11 and X30 and X71) xor (X11 and X30 and X73) xor (X11 and X31 and X73) xor (X11 and X33 and X70) xor (X11 and X33 and X71) xor (X11 and X33 and X73) xor (X13 and X30 and X71) xor (X13 and X31 and X70) xor (X13 and X31 and X71) xor (X13 and X31 and X73) xor (X13 and X33 and X70) xor (X20 and X30 and X71) xor (X20 and X31 and X70) xor (X20 and X31 and X73) xor (X20 and X33 and X71) xor (X20 and X33 and X73) xor (X21 and X30 and X71) xor (X21 and X30 and X73) xor (X21 and X31 and X73) xor (X21 and X33 and X70) xor (X21 and X33 and X71) xor (X21 and X33 and X73) xor (X23 and X30 and X71) xor (X23 and X31 and X70) xor (X23 and X31 and X71) xor (X23 and X31 and X73) xor (X23 and X33 and X70) xor (X20 and X40 and X71) xor (X20 and X41 and X70) xor (X20 and X41 and X73) xor (X20 and X43 and X71) xor (X20 and X43 and X73) xor (X21 and X40 and X71) xor (X21 and X40 and X73) xor (X21 and X41 and X73) xor (X21 and X43 and X70) xor (X21 and X43 and X71) xor (X21 and X43 and X73) xor (X23 and X40 and X71) xor (X23 and X41 and X70) xor (X23 and X41 and X71) xor (X23 and X41 and X73) xor (X23 and X43 and X70) xor (X20 and X50 and X71) xor (X20 and X51 and X70) xor (X20 and X51 and X73) xor (X20 and X53 and X71) xor (X20 and X53 and X73) xor (X21 and X50 and X71) xor (X21 and X50 and X73) xor (X21 and X51 and X73) xor (X21 and X53 and X70) xor (X21 and X53 and X71) xor (X21 and X53 and X73) xor (X23 and X50 and X71) xor (X23 and X51 and X70) xor (X23 and X51 and X71) xor (X23 and X51 and X73) xor (X23 and X53 and X70) xor (X10 and X60 and X71) xor (X10 and X61 and X70) xor (X10 and X61 and X73) xor (X10 and X63 and X71) xor (X10 and X63 and X73) xor (X11 and X60 and X71) xor (X11 and X60 and X73) xor (X11 and X61 and X73) xor (X11 and X63 and X70) xor (X11 and X63 and X71) xor (X11 and X63 and X73) xor (X13 and X60 and X71) xor (X13 and X61 and X70) xor (X13 and X61 and X71) xor (X13 and X61 and X73) xor (X13 and X63 and X70) xor (X20 and X60 and X71) xor (X20 and X61 and X70) xor (X20 and X61 and X73) xor (X20 and X63 and X71) xor (X20 and X63 and X73) xor (X21 and X60 and X71) xor (X21 and X60 and X73) xor (X21 and X61 and X73) xor (X21 and X63 and X70) xor (X21 and X63 and X71) xor (X21 and X63 and X73) xor (X23 and X60 and X71) xor (X23 and X61 and X70) xor (X23 and X61 and X71) xor (X23 and X61 and X73) xor (X23 and X63 and X70) xor (X40 and X60 and X71) xor (X40 and X61 and X70) xor (X40 and X61 and X73) xor (X40 and X63 and X71) xor (X40 and X63 and X73) xor (X41 and X60 and X71) xor (X41 and X60 and X73) xor (X41 and X61 and X73) xor (X41 and X63 and X70) xor (X41 and X63 and X71) xor (X41 and X63 and X73) xor (X43 and X60 and X71) xor (X43 and X61 and X70) xor (X43 and X61 and X71) xor (X43 and X61 and X73) xor (X43 and X63 and X70) xor (X50 and X60 and X71) xor (X50 and X61 and X70) xor (X50 and X61 and X73) xor (X50 and X63 and X71) xor (X50 and X63 and X73) xor (X51 and X60 and X71) xor (X51 and X60 and X73) xor (X51 and X61 and X73) xor (X51 and X63 and X70) xor (X51 and X63 and X71) xor (X51 and X63 and X73) xor (X53 and X60 and X71) xor (X53 and X61 and X70) xor (X53 and X61 and X71) xor (X53 and X61 and X73) xor (X53 and X63 and X70));
    F20  <= ((X00 and X10) xor (X00 and X11) xor (X02 and X10) xor (X00 and X12) xor (X20) xor (X30) xor (X10 and X30) xor (X10 and X31) xor (X12 and X30) xor (X10 and X32) xor (X10 and X20 and X30) xor (X10 and X20 and X32) xor (X10 and X21 and X31) xor (X10 and X21 and X32) xor (X10 and X22 and X31) xor (X11 and X20 and X30) xor (X11 and X20 and X32) xor (X11 and X21 and X30) xor (X11 and X22 and X30) xor (X11 and X22 and X31) xor (X12 and X20 and X30) xor (X12 and X20 and X31) xor (X12 and X21 and X30) xor (X12 and X21 and X31) xor (X12 and X22 and X30) xor (X12 and X22 and X32) xor (X40) xor (X00 and X20 and X40) xor (X00 and X20 and X42) xor (X00 and X21 and X41) xor (X00 and X21 and X42) xor (X00 and X22 and X41) xor (X0_1 and X20 and X40) xor (X0_1 and X20 and X42) xor (X0_1 and X21 and X40) xor (X0_1 and X22 and X40) xor (X0_1 and X22 and X41) xor (X02 and X20 and X40) xor (X02 and X20 and X41) xor (X02 and X21 and X40) xor (X02 and X21 and X41) xor (X02 and X22 and X40) xor (X02 and X22 and X42) xor (X10 and X20 and X40) xor (X10 and X20 and X42) xor (X10 and X21 and X41) xor (X10 and X21 and X42) xor (X10 and X22 and X41) xor (X11 and X20 and X40) xor (X11 and X20 and X42) xor (X11 and X21 and X40) xor (X11 and X22 and X40) xor (X11 and X22 and X41) xor (X12 and X20 and X40) xor (X12 and X20 and X41) xor (X12 and X21 and X40) xor (X12 and X21 and X41) xor (X12 and X22 and X40) xor (X12 and X22 and X42) xor (X30 and X40) xor (X30 and X41) xor (X32 and X40) xor (X30 and X42) xor (X10 and X30 and X40) xor (X10 and X30 and X42) xor (X10 and X31 and X41) xor (X10 and X31 and X42) xor (X10 and X32 and X41) xor (X11 and X30 and X40) xor (X11 and X30 and X42) xor (X11 and X31 and X40) xor (X11 and X32 and X40) xor (X11 and X32 and X41) xor (X12 and X30 and X40) xor (X12 and X30 and X41) xor (X12 and X31 and X40) xor (X12 and X31 and X41) xor (X12 and X32 and X40) xor (X12 and X32 and X42) xor (X20 and X30 and X40) xor (X20 and X30 and X42) xor (X20 and X31 and X41) xor (X20 and X31 and X42) xor (X20 and X32 and X41) xor (X21 and X30 and X40) xor (X21 and X30 and X42) xor (X21 and X31 and X40) xor (X21 and X32 and X40) xor (X21 and X32 and X41) xor (X22 and X30 and X40) xor (X22 and X30 and X41) xor (X22 and X31 and X40) xor (X22 and X31 and X41) xor (X22 and X32 and X40) xor (X22 and X32 and X42) xor (X00 and X50) xor (X00 and X51) xor (X02 and X50) xor (X00 and X52) xor (X20 and X50) xor (X20 and X51) xor (X22 and X50) xor (X20 and X52) xor (X00 and X20 and X50) xor (X00 and X20 and X52) xor (X00 and X21 and X51) xor (X00 and X21 and X52) xor (X00 and X22 and X51) xor (X0_1 and X20 and X50) xor (X0_1 and X20 and X52) xor (X0_1 and X21 and X50) xor (X0_1 and X22 and X50) xor (X0_1 and X22 and X51) xor (X02 and X20 and X50) xor (X02 and X20 and X51) xor (X02 and X21 and X50) xor (X02 and X21 and X51) xor (X02 and X22 and X50) xor (X02 and X22 and X52) xor (X30 and X50) xor (X30 and X51) xor (X32 and X50) xor (X30 and X52) xor (X00 and X30 and X50) xor (X00 and X30 and X52) xor (X00 and X31 and X51) xor (X00 and X31 and X52) xor (X00 and X32 and X51) xor (X0_1 and X30 and X50) xor (X0_1 and X30 and X52) xor (X0_1 and X31 and X50) xor (X0_1 and X32 and X50) xor (X0_1 and X32 and X51) xor (X02 and X30 and X50) xor (X02 and X30 and X51) xor (X02 and X31 and X50) xor (X02 and X31 and X51) xor (X02 and X32 and X50) xor (X02 and X32 and X52) xor (X10 and X30 and X50) xor (X10 and X30 and X52) xor (X10 and X31 and X51) xor (X10 and X31 and X52) xor (X10 and X32 and X51) xor (X11 and X30 and X50) xor (X11 and X30 and X52) xor (X11 and X31 and X50) xor (X11 and X32 and X50) xor (X11 and X32 and X51) xor (X12 and X30 and X50) xor (X12 and X30 and X51) xor (X12 and X31 and X50) xor (X12 and X31 and X51) xor (X12 and X32 and X50) xor (X12 and X32 and X52) xor (X40 and X50) xor (X40 and X51) xor (X42 and X50) xor (X40 and X52) xor (X00 and X40 and X50) xor (X00 and X40 and X52) xor (X00 and X41 and X51) xor (X00 and X41 and X52) xor (X00 and X42 and X51) xor (X0_1 and X40 and X50) xor (X0_1 and X40 and X52) xor (X0_1 and X41 and X50) xor (X0_1 and X42 and X50) xor (X0_1 and X42 and X51) xor (X02 and X40 and X50) xor (X02 and X40 and X51) xor (X02 and X41 and X50) xor (X02 and X41 and X51) xor (X02 and X42 and X50) xor (X02 and X42 and X52) xor (X20 and X40 and X50) xor (X20 and X40 and X52) xor (X20 and X41 and X51) xor (X20 and X41 and X52) xor (X20 and X42 and X51) xor (X21 and X40 and X50) xor (X21 and X40 and X52) xor (X21 and X41 and X50) xor (X21 and X42 and X50) xor (X21 and X42 and X51) xor (X22 and X40 and X50) xor (X22 and X40 and X51) xor (X22 and X41 and X50) xor (X22 and X41 and X51) xor (X22 and X42 and X50) xor (X22 and X42 and X52) xor (X30 and X40 and X50) xor (X30 and X40 and X52) xor (X30 and X41 and X51) xor (X30 and X41 and X52) xor (X30 and X42 and X51) xor (X31 and X40 and X50) xor (X31 and X40 and X52) xor (X31 and X41 and X50) xor (X31 and X42 and X50) xor (X31 and X42 and X51) xor (X32 and X40 and X50) xor (X32 and X40 and X51) xor (X32 and X41 and X50) xor (X32 and X41 and X51) xor (X32 and X42 and X50) xor (X32 and X42 and X52) xor (X10 and X20 and X60) xor (X10 and X20 and X62) xor (X10 and X21 and X61) xor (X10 and X21 and X62) xor (X10 and X22 and X61) xor (X11 and X20 and X60) xor (X11 and X20 and X62) xor (X11 and X21 and X60) xor (X11 and X22 and X60) xor (X11 and X22 and X61) xor (X12 and X20 and X60) xor (X12 and X20 and X61) xor (X12 and X21 and X60) xor (X12 and X21 and X61) xor (X12 and X22 and X60) xor (X12 and X22 and X62) xor (X30 and X60) xor (X30 and X61) xor (X32 and X60) xor (X30 and X62) xor (X00 and X30 and X60) xor (X00 and X30 and X62) xor (X00 and X31 and X61) xor (X00 and X31 and X62) xor (X00 and X32 and X61) xor (X0_1 and X30 and X60) xor (X0_1 and X30 and X62) xor (X0_1 and X31 and X60) xor (X0_1 and X32 and X60) xor (X0_1 and X32 and X61) xor (X02 and X30 and X60) xor (X02 and X30 and X61) xor (X02 and X31 and X60) xor (X02 and X31 and X61) xor (X02 and X32 and X60) xor (X02 and X32 and X62) xor (X10 and X30 and X60) xor (X10 and X30 and X62) xor (X10 and X31 and X61) xor (X10 and X31 and X62) xor (X10 and X32 and X61) xor (X11 and X30 and X60) xor (X11 and X30 and X62) xor (X11 and X31 and X60) xor (X11 and X32 and X60) xor (X11 and X32 and X61) xor (X12 and X30 and X60) xor (X12 and X30 and X61) xor (X12 and X31 and X60) xor (X12 and X31 and X61) xor (X12 and X32 and X60) xor (X12 and X32 and X62) xor (X20 and X30 and X60) xor (X20 and X30 and X62) xor (X20 and X31 and X61) xor (X20 and X31 and X62) xor (X20 and X32 and X61) xor (X21 and X30 and X60) xor (X21 and X30 and X62) xor (X21 and X31 and X60) xor (X21 and X32 and X60) xor (X21 and X32 and X61) xor (X22 and X30 and X60) xor (X22 and X30 and X61) xor (X22 and X31 and X60) xor (X22 and X31 and X61) xor (X22 and X32 and X60) xor (X22 and X32 and X62) xor (X50 and X60) xor (X50 and X61) xor (X52 and X60) xor (X50 and X62) xor (X00 and X50 and X60) xor (X00 and X50 and X62) xor (X00 and X51 and X61) xor (X00 and X51 and X62) xor (X00 and X52 and X61) xor (X0_1 and X50 and X60) xor (X0_1 and X50 and X62) xor (X0_1 and X51 and X60) xor (X0_1 and X52 and X60) xor (X0_1 and X52 and X61) xor (X02 and X50 and X60) xor (X02 and X50 and X61) xor (X02 and X51 and X60) xor (X02 and X51 and X61) xor (X02 and X52 and X60) xor (X02 and X52 and X62) xor (X10 and X50 and X60) xor (X10 and X50 and X62) xor (X10 and X51 and X61) xor (X10 and X51 and X62) xor (X10 and X52 and X61) xor (X11 and X50 and X60) xor (X11 and X50 and X62) xor (X11 and X51 and X60) xor (X11 and X52 and X60) xor (X11 and X52 and X61) xor (X12 and X50 and X60) xor (X12 and X50 and X61) xor (X12 and X51 and X60) xor (X12 and X51 and X61) xor (X12 and X52 and X60) xor (X12 and X52 and X62) xor (X20 and X50 and X60) xor (X20 and X50 and X62) xor (X20 and X51 and X61) xor (X20 and X51 and X62) xor (X20 and X52 and X61) xor (X21 and X50 and X60) xor (X21 and X50 and X62) xor (X21 and X51 and X60) xor (X21 and X52 and X60) xor (X21 and X52 and X61) xor (X22 and X50 and X60) xor (X22 and X50 and X61) xor (X22 and X51 and X60) xor (X22 and X51 and X61) xor (X22 and X52 and X60) xor (X22 and X52 and X62) xor (X40 and X50 and X60) xor (X40 and X50 and X62) xor (X40 and X51 and X61) xor (X40 and X51 and X62) xor (X40 and X52 and X61) xor (X41 and X50 and X60) xor (X41 and X50 and X62) xor (X41 and X51 and X60) xor (X41 and X52 and X60) xor (X41 and X52 and X61) xor (X42 and X50 and X60) xor (X42 and X50 and X61) xor (X42 and X51 and X60) xor (X42 and X51 and X61) xor (X42 and X52 and X60) xor (X42 and X52 and X62) xor (X70) xor (X10 and X70) xor (X10 and X71) xor (X12 and X70) xor (X10 and X72) xor (X00 and X10 and X70) xor (X00 and X10 and X72) xor (X00 and X11 and X71) xor (X00 and X11 and X72) xor (X00 and X12 and X71) xor (X0_1 and X10 and X70) xor (X0_1 and X10 and X72) xor (X0_1 and X11 and X70) xor (X0_1 and X12 and X70) xor (X0_1 and X12 and X71) xor (X02 and X10 and X70) xor (X02 and X10 and X71) xor (X02 and X11 and X70) xor (X02 and X11 and X71) xor (X02 and X12 and X70) xor (X02 and X12 and X72) xor (X10 and X20 and X70) xor (X10 and X20 and X72) xor (X10 and X21 and X71) xor (X10 and X21 and X72) xor (X10 and X22 and X71) xor (X11 and X20 and X70) xor (X11 and X20 and X72) xor (X11 and X21 and X70) xor (X11 and X22 and X70) xor (X11 and X22 and X71) xor (X12 and X20 and X70) xor (X12 and X20 and X71) xor (X12 and X21 and X70) xor (X12 and X21 and X71) xor (X12 and X22 and X70) xor (X12 and X22 and X72) xor (X30 and X70) xor (X30 and X71) xor (X32 and X70) xor (X30 and X72) xor (X00 and X30 and X70) xor (X00 and X30 and X72) xor (X00 and X31 and X71) xor (X00 and X31 and X72) xor (X00 and X32 and X71) xor (X0_1 and X30 and X70) xor (X0_1 and X30 and X72) xor (X0_1 and X31 and X70) xor (X0_1 and X32 and X70) xor (X0_1 and X32 and X71) xor (X02 and X30 and X70) xor (X02 and X30 and X71) xor (X02 and X31 and X70) xor (X02 and X31 and X71) xor (X02 and X32 and X70) xor (X02 and X32 and X72) xor (X40 and X70) xor (X40 and X71) xor (X42 and X70) xor (X40 and X72) xor (X00 and X40 and X70) xor (X00 and X40 and X72) xor (X00 and X41 and X71) xor (X00 and X41 and X72) xor (X00 and X42 and X71) xor (X0_1 and X40 and X70) xor (X0_1 and X40 and X72) xor (X0_1 and X41 and X70) xor (X0_1 and X42 and X70) xor (X0_1 and X42 and X71) xor (X02 and X40 and X70) xor (X02 and X40 and X71) xor (X02 and X41 and X70) xor (X02 and X41 and X71) xor (X02 and X42 and X70) xor (X02 and X42 and X72) xor (X10 and X40 and X70) xor (X10 and X40 and X72) xor (X10 and X41 and X71) xor (X10 and X41 and X72) xor (X10 and X42 and X71) xor (X11 and X40 and X70) xor (X11 and X40 and X72) xor (X11 and X41 and X70) xor (X11 and X42 and X70) xor (X11 and X42 and X71) xor (X12 and X40 and X70) xor (X12 and X40 and X71) xor (X12 and X41 and X70) xor (X12 and X41 and X71) xor (X12 and X42 and X70) xor (X12 and X42 and X72) xor (X30 and X40 and X70) xor (X30 and X40 and X72) xor (X30 and X41 and X71) xor (X30 and X41 and X72) xor (X30 and X42 and X71) xor (X31 and X40 and X70) xor (X31 and X40 and X72) xor (X31 and X41 and X70) xor (X31 and X42 and X70) xor (X31 and X42 and X71) xor (X32 and X40 and X70) xor (X32 and X40 and X71) xor (X32 and X41 and X70) xor (X32 and X41 and X71) xor (X32 and X42 and X70) xor (X32 and X42 and X72) xor (X50 and X70) xor (X50 and X71) xor (X52 and X70) xor (X50 and X72) xor (X00 and X50 and X70) xor (X00 and X50 and X72) xor (X00 and X51 and X71) xor (X00 and X51 and X72) xor (X00 and X52 and X71) xor (X0_1 and X50 and X70) xor (X0_1 and X50 and X72) xor (X0_1 and X51 and X70) xor (X0_1 and X52 and X70) xor (X0_1 and X52 and X71) xor (X02 and X50 and X70) xor (X02 and X50 and X71) xor (X02 and X51 and X70) xor (X02 and X51 and X71) xor (X02 and X52 and X70) xor (X02 and X52 and X72) xor (X10 and X50 and X70) xor (X10 and X50 and X72) xor (X10 and X51 and X71) xor (X10 and X51 and X72) xor (X10 and X52 and X71) xor (X11 and X50 and X70) xor (X11 and X50 and X72) xor (X11 and X51 and X70) xor (X11 and X52 and X70) xor (X11 and X52 and X71) xor (X12 and X50 and X70) xor (X12 and X50 and X71) xor (X12 and X51 and X70) xor (X12 and X51 and X71) xor (X12 and X52 and X70) xor (X12 and X52 and X72) xor (X60 and X70) xor (X60 and X71) xor (X62 and X70) xor (X60 and X72) xor (X00 and X60 and X70) xor (X00 and X60 and X72) xor (X00 and X61 and X71) xor (X00 and X61 and X72) xor (X00 and X62 and X71) xor (X0_1 and X60 and X70) xor (X0_1 and X60 and X72) xor (X0_1 and X61 and X70) xor (X0_1 and X62 and X70) xor (X0_1 and X62 and X71) xor (X02 and X60 and X70) xor (X02 and X60 and X71) xor (X02 and X61 and X70) xor (X02 and X61 and X71) xor (X02 and X62 and X70) xor (X02 and X62 and X72) xor (X10 and X60 and X70) xor (X10 and X60 and X72) xor (X10 and X61 and X71) xor (X10 and X61 and X72) xor (X10 and X62 and X71) xor (X11 and X60 and X70) xor (X11 and X60 and X72) xor (X11 and X61 and X70) xor (X11 and X62 and X70) xor (X11 and X62 and X71) xor (X12 and X60 and X70) xor (X12 and X60 and X71) xor (X12 and X61 and X70) xor (X12 and X61 and X71) xor (X12 and X62 and X70) xor (X12 and X62 and X72) xor (X40 and X60 and X70) xor (X40 and X60 and X72) xor (X40 and X61 and X71) xor (X40 and X61 and X72) xor (X40 and X62 and X71) xor (X41 and X60 and X70) xor (X41 and X60 and X72) xor (X41 and X61 and X70) xor (X41 and X62 and X70) xor (X41 and X62 and X71) xor (X42 and X60 and X70) xor (X42 and X60 and X71) xor (X42 and X61 and X70) xor (X42 and X61 and X71) xor (X42 and X62 and X70) xor (X42 and X62 and X72));
    F21  <= ((X0_1 and X11) xor (X0_1 and X12) xor (X02 and X11) xor (X0_1 and X13) xor (X21) xor (X31) xor (X11 and X31) xor (X11 and X32) xor (X12 and X31) xor (X11 and X33) xor (X11 and X21 and X31) xor (X11 and X21 and X32) xor (X11 and X22 and X32) xor (X11 and X22 and X33) xor (X11 and X23 and X32) xor (X12 and X21 and X32) xor (X12 and X21 and X33) xor (X12 and X22 and X31) xor (X12 and X22 and X33) xor (X12 and X23 and X31) xor (X12 and X23 and X32) xor (X13 and X21 and X32) xor (X13 and X22 and X31) xor (X13 and X22 and X33) xor (X13 and X23 and X31) xor (X13 and X23 and X33) xor (X41) xor (X0_1 and X21 and X41) xor (X0_1 and X21 and X42) xor (X0_1 and X22 and X42) xor (X0_1 and X22 and X43) xor (X0_1 and X23 and X42) xor (X02 and X21 and X42) xor (X02 and X21 and X43) xor (X02 and X22 and X41) xor (X02 and X22 and X43) xor (X02 and X23 and X41) xor (X02 and X23 and X42) xor (X03 and X21 and X42) xor (X03 and X22 and X41) xor (X03 and X22 and X43) xor (X03 and X23 and X41) xor (X03 and X23 and X43) xor (X11 and X21 and X41) xor (X11 and X21 and X42) xor (X11 and X22 and X42) xor (X11 and X22 and X43) xor (X11 and X23 and X42) xor (X12 and X21 and X42) xor (X12 and X21 and X43) xor (X12 and X22 and X41) xor (X12 and X22 and X43) xor (X12 and X23 and X41) xor (X12 and X23 and X42) xor (X13 and X21 and X42) xor (X13 and X22 and X41) xor (X13 and X22 and X43) xor (X13 and X23 and X41) xor (X13 and X23 and X43) xor (X31 and X41) xor (X31 and X42) xor (X32 and X41) xor (X31 and X43) xor (X11 and X31 and X41) xor (X11 and X31 and X42) xor (X11 and X32 and X42) xor (X11 and X32 and X43) xor (X11 and X33 and X42) xor (X12 and X31 and X42) xor (X12 and X31 and X43) xor (X12 and X32 and X41) xor (X12 and X32 and X43) xor (X12 and X33 and X41) xor (X12 and X33 and X42) xor (X13 and X31 and X42) xor (X13 and X32 and X41) xor (X13 and X32 and X43) xor (X13 and X33 and X41) xor (X13 and X33 and X43) xor (X21 and X31 and X41) xor (X21 and X31 and X42) xor (X21 and X32 and X42) xor (X21 and X32 and X43) xor (X21 and X33 and X42) xor (X22 and X31 and X42) xor (X22 and X31 and X43) xor (X22 and X32 and X41) xor (X22 and X32 and X43) xor (X22 and X33 and X41) xor (X22 and X33 and X42) xor (X23 and X31 and X42) xor (X23 and X32 and X41) xor (X23 and X32 and X43) xor (X23 and X33 and X41) xor (X23 and X33 and X43) xor (X0_1 and X51) xor (X0_1 and X52) xor (X02 and X51) xor (X0_1 and X53) xor (X21 and X51) xor (X21 and X52) xor (X22 and X51) xor (X21 and X53) xor (X0_1 and X21 and X51) xor (X0_1 and X21 and X52) xor (X0_1 and X22 and X52) xor (X0_1 and X22 and X53) xor (X0_1 and X23 and X52) xor (X02 and X21 and X52) xor (X02 and X21 and X53) xor (X02 and X22 and X51) xor (X02 and X22 and X53) xor (X02 and X23 and X51) xor (X02 and X23 and X52) xor (X03 and X21 and X52) xor (X03 and X22 and X51) xor (X03 and X22 and X53) xor (X03 and X23 and X51) xor (X03 and X23 and X53) xor (X31 and X51) xor (X31 and X52) xor (X32 and X51) xor (X31 and X53) xor (X0_1 and X31 and X51) xor (X0_1 and X31 and X52) xor (X0_1 and X32 and X52) xor (X0_1 and X32 and X53) xor (X0_1 and X33 and X52) xor (X02 and X31 and X52) xor (X02 and X31 and X53) xor (X02 and X32 and X51) xor (X02 and X32 and X53) xor (X02 and X33 and X51) xor (X02 and X33 and X52) xor (X03 and X31 and X52) xor (X03 and X32 and X51) xor (X03 and X32 and X53) xor (X03 and X33 and X51) xor (X03 and X33 and X53) xor (X11 and X31 and X51) xor (X11 and X31 and X52) xor (X11 and X32 and X52) xor (X11 and X32 and X53) xor (X11 and X33 and X52) xor (X12 and X31 and X52) xor (X12 and X31 and X53) xor (X12 and X32 and X51) xor (X12 and X32 and X53) xor (X12 and X33 and X51) xor (X12 and X33 and X52) xor (X13 and X31 and X52) xor (X13 and X32 and X51) xor (X13 and X32 and X53) xor (X13 and X33 and X51) xor (X13 and X33 and X53) xor (X41 and X51) xor (X41 and X52) xor (X42 and X51) xor (X41 and X53) xor (X0_1 and X41 and X51) xor (X0_1 and X41 and X52) xor (X0_1 and X42 and X52) xor (X0_1 and X42 and X53) xor (X0_1 and X43 and X52) xor (X02 and X41 and X52) xor (X02 and X41 and X53) xor (X02 and X42 and X51) xor (X02 and X42 and X53) xor (X02 and X43 and X51) xor (X02 and X43 and X52) xor (X03 and X41 and X52) xor (X03 and X42 and X51) xor (X03 and X42 and X53) xor (X03 and X43 and X51) xor (X03 and X43 and X53) xor (X21 and X41 and X51) xor (X21 and X41 and X52) xor (X21 and X42 and X52) xor (X21 and X42 and X53) xor (X21 and X43 and X52) xor (X22 and X41 and X52) xor (X22 and X41 and X53) xor (X22 and X42 and X51) xor (X22 and X42 and X53) xor (X22 and X43 and X51) xor (X22 and X43 and X52) xor (X23 and X41 and X52) xor (X23 and X42 and X51) xor (X23 and X42 and X53) xor (X23 and X43 and X51) xor (X23 and X43 and X53) xor (X31 and X41 and X51) xor (X31 and X41 and X52) xor (X31 and X42 and X52) xor (X31 and X42 and X53) xor (X31 and X43 and X52) xor (X32 and X41 and X52) xor (X32 and X41 and X53) xor (X32 and X42 and X51) xor (X32 and X42 and X53) xor (X32 and X43 and X51) xor (X32 and X43 and X52) xor (X33 and X41 and X52) xor (X33 and X42 and X51) xor (X33 and X42 and X53) xor (X33 and X43 and X51) xor (X33 and X43 and X53) xor (X11 and X21 and X61) xor (X11 and X21 and X62) xor (X11 and X22 and X62) xor (X11 and X22 and X63) xor (X11 and X23 and X62) xor (X12 and X21 and X62) xor (X12 and X21 and X63) xor (X12 and X22 and X61) xor (X12 and X22 and X63) xor (X12 and X23 and X61) xor (X12 and X23 and X62) xor (X13 and X21 and X62) xor (X13 and X22 and X61) xor (X13 and X22 and X63) xor (X13 and X23 and X61) xor (X13 and X23 and X63) xor (X31 and X61) xor (X31 and X62) xor (X32 and X61) xor (X31 and X63) xor (X0_1 and X31 and X61) xor (X0_1 and X31 and X62) xor (X0_1 and X32 and X62) xor (X0_1 and X32 and X63) xor (X0_1 and X33 and X62) xor (X02 and X31 and X62) xor (X02 and X31 and X63) xor (X02 and X32 and X61) xor (X02 and X32 and X63) xor (X02 and X33 and X61) xor (X02 and X33 and X62) xor (X03 and X31 and X62) xor (X03 and X32 and X61) xor (X03 and X32 and X63) xor (X03 and X33 and X61) xor (X03 and X33 and X63) xor (X11 and X31 and X61) xor (X11 and X31 and X62) xor (X11 and X32 and X62) xor (X11 and X32 and X63) xor (X11 and X33 and X62) xor (X12 and X31 and X62) xor (X12 and X31 and X63) xor (X12 and X32 and X61) xor (X12 and X32 and X63) xor (X12 and X33 and X61) xor (X12 and X33 and X62) xor (X13 and X31 and X62) xor (X13 and X32 and X61) xor (X13 and X32 and X63) xor (X13 and X33 and X61) xor (X13 and X33 and X63) xor (X21 and X31 and X61) xor (X21 and X31 and X62) xor (X21 and X32 and X62) xor (X21 and X32 and X63) xor (X21 and X33 and X62) xor (X22 and X31 and X62) xor (X22 and X31 and X63) xor (X22 and X32 and X61) xor (X22 and X32 and X63) xor (X22 and X33 and X61) xor (X22 and X33 and X62) xor (X23 and X31 and X62) xor (X23 and X32 and X61) xor (X23 and X32 and X63) xor (X23 and X33 and X61) xor (X23 and X33 and X63) xor (X51 and X61) xor (X51 and X62) xor (X52 and X61) xor (X51 and X63) xor (X0_1 and X51 and X61) xor (X0_1 and X51 and X62) xor (X0_1 and X52 and X62) xor (X0_1 and X52 and X63) xor (X0_1 and X53 and X62) xor (X02 and X51 and X62) xor (X02 and X51 and X63) xor (X02 and X52 and X61) xor (X02 and X52 and X63) xor (X02 and X53 and X61) xor (X02 and X53 and X62) xor (X03 and X51 and X62) xor (X03 and X52 and X61) xor (X03 and X52 and X63) xor (X03 and X53 and X61) xor (X03 and X53 and X63) xor (X11 and X51 and X61) xor (X11 and X51 and X62) xor (X11 and X52 and X62) xor (X11 and X52 and X63) xor (X11 and X53 and X62) xor (X12 and X51 and X62) xor (X12 and X51 and X63) xor (X12 and X52 and X61) xor (X12 and X52 and X63) xor (X12 and X53 and X61) xor (X12 and X53 and X62) xor (X13 and X51 and X62) xor (X13 and X52 and X61) xor (X13 and X52 and X63) xor (X13 and X53 and X61) xor (X13 and X53 and X63) xor (X21 and X51 and X61) xor (X21 and X51 and X62) xor (X21 and X52 and X62) xor (X21 and X52 and X63) xor (X21 and X53 and X62) xor (X22 and X51 and X62) xor (X22 and X51 and X63) xor (X22 and X52 and X61) xor (X22 and X52 and X63) xor (X22 and X53 and X61) xor (X22 and X53 and X62) xor (X23 and X51 and X62) xor (X23 and X52 and X61) xor (X23 and X52 and X63) xor (X23 and X53 and X61) xor (X23 and X53 and X63) xor (X41 and X51 and X61) xor (X41 and X51 and X62) xor (X41 and X52 and X62) xor (X41 and X52 and X63) xor (X41 and X53 and X62) xor (X42 and X51 and X62) xor (X42 and X51 and X63) xor (X42 and X52 and X61) xor (X42 and X52 and X63) xor (X42 and X53 and X61) xor (X42 and X53 and X62) xor (X43 and X51 and X62) xor (X43 and X52 and X61) xor (X43 and X52 and X63) xor (X43 and X53 and X61) xor (X43 and X53 and X63) xor (X71) xor (X11 and X71) xor (X11 and X72) xor (X12 and X71) xor (X11 and X73) xor (X0_1 and X11 and X71) xor (X0_1 and X11 and X72) xor (X0_1 and X12 and X72) xor (X0_1 and X12 and X73) xor (X0_1 and X13 and X72) xor (X02 and X11 and X72) xor (X02 and X11 and X73) xor (X02 and X12 and X71) xor (X02 and X12 and X73) xor (X02 and X13 and X71) xor (X02 and X13 and X72) xor (X03 and X11 and X72) xor (X03 and X12 and X71) xor (X03 and X12 and X73) xor (X03 and X13 and X71) xor (X03 and X13 and X73) xor (X11 and X21 and X71) xor (X11 and X21 and X72) xor (X11 and X22 and X72) xor (X11 and X22 and X73) xor (X11 and X23 and X72) xor (X12 and X21 and X72) xor (X12 and X21 and X73) xor (X12 and X22 and X71) xor (X12 and X22 and X73) xor (X12 and X23 and X71) xor (X12 and X23 and X72) xor (X13 and X21 and X72) xor (X13 and X22 and X71) xor (X13 and X22 and X73) xor (X13 and X23 and X71) xor (X13 and X23 and X73) xor (X31 and X71) xor (X31 and X72) xor (X32 and X71) xor (X31 and X73) xor (X0_1 and X31 and X71) xor (X0_1 and X31 and X72) xor (X0_1 and X32 and X72) xor (X0_1 and X32 and X73) xor (X0_1 and X33 and X72) xor (X02 and X31 and X72) xor (X02 and X31 and X73) xor (X02 and X32 and X71) xor (X02 and X32 and X73) xor (X02 and X33 and X71) xor (X02 and X33 and X72) xor (X03 and X31 and X72) xor (X03 and X32 and X71) xor (X03 and X32 and X73) xor (X03 and X33 and X71) xor (X03 and X33 and X73) xor (X41 and X71) xor (X41 and X72) xor (X42 and X71) xor (X41 and X73) xor (X0_1 and X41 and X71) xor (X0_1 and X41 and X72) xor (X0_1 and X42 and X72) xor (X0_1 and X42 and X73) xor (X0_1 and X43 and X72) xor (X02 and X41 and X72) xor (X02 and X41 and X73) xor (X02 and X42 and X71) xor (X02 and X42 and X73) xor (X02 and X43 and X71) xor (X02 and X43 and X72) xor (X03 and X41 and X72) xor (X03 and X42 and X71) xor (X03 and X42 and X73) xor (X03 and X43 and X71) xor (X03 and X43 and X73) xor (X11 and X41 and X71) xor (X11 and X41 and X72) xor (X11 and X42 and X72) xor (X11 and X42 and X73) xor (X11 and X43 and X72) xor (X12 and X41 and X72) xor (X12 and X41 and X73) xor (X12 and X42 and X71) xor (X12 and X42 and X73) xor (X12 and X43 and X71) xor (X12 and X43 and X72) xor (X13 and X41 and X72) xor (X13 and X42 and X71) xor (X13 and X42 and X73) xor (X13 and X43 and X71) xor (X13 and X43 and X73) xor (X31 and X41 and X71) xor (X31 and X41 and X72) xor (X31 and X42 and X72) xor (X31 and X42 and X73) xor (X31 and X43 and X72) xor (X32 and X41 and X72) xor (X32 and X41 and X73) xor (X32 and X42 and X71) xor (X32 and X42 and X73) xor (X32 and X43 and X71) xor (X32 and X43 and X72) xor (X33 and X41 and X72) xor (X33 and X42 and X71) xor (X33 and X42 and X73) xor (X33 and X43 and X71) xor (X33 and X43 and X73) xor (X51 and X71) xor (X51 and X72) xor (X52 and X71) xor (X51 and X73) xor (X0_1 and X51 and X71) xor (X0_1 and X51 and X72) xor (X0_1 and X52 and X72) xor (X0_1 and X52 and X73) xor (X0_1 and X53 and X72) xor (X02 and X51 and X72) xor (X02 and X51 and X73) xor (X02 and X52 and X71) xor (X02 and X52 and X73) xor (X02 and X53 and X71) xor (X02 and X53 and X72) xor (X03 and X51 and X72) xor (X03 and X52 and X71) xor (X03 and X52 and X73) xor (X03 and X53 and X71) xor (X03 and X53 and X73) xor (X11 and X51 and X71) xor (X11 and X51 and X72) xor (X11 and X52 and X72) xor (X11 and X52 and X73) xor (X11 and X53 and X72) xor (X12 and X51 and X72) xor (X12 and X51 and X73) xor (X12 and X52 and X71) xor (X12 and X52 and X73) xor (X12 and X53 and X71) xor (X12 and X53 and X72) xor (X13 and X51 and X72) xor (X13 and X52 and X71) xor (X13 and X52 and X73) xor (X13 and X53 and X71) xor (X13 and X53 and X73) xor (X61 and X71) xor (X61 and X72) xor (X62 and X71) xor (X61 and X73) xor (X0_1 and X61 and X71) xor (X0_1 and X61 and X72) xor (X0_1 and X62 and X72) xor (X0_1 and X62 and X73) xor (X0_1 and X63 and X72) xor (X02 and X61 and X72) xor (X02 and X61 and X73) xor (X02 and X62 and X71) xor (X02 and X62 and X73) xor (X02 and X63 and X71) xor (X02 and X63 and X72) xor (X03 and X61 and X72) xor (X03 and X62 and X71) xor (X03 and X62 and X73) xor (X03 and X63 and X71) xor (X03 and X63 and X73) xor (X11 and X61 and X71) xor (X11 and X61 and X72) xor (X11 and X62 and X72) xor (X11 and X62 and X73) xor (X11 and X63 and X72) xor (X12 and X61 and X72) xor (X12 and X61 and X73) xor (X12 and X62 and X71) xor (X12 and X62 and X73) xor (X12 and X63 and X71) xor (X12 and X63 and X72) xor (X13 and X61 and X72) xor (X13 and X62 and X71) xor (X13 and X62 and X73) xor (X13 and X63 and X71) xor (X13 and X63 and X73) xor (X41 and X61 and X71) xor (X41 and X61 and X72) xor (X41 and X62 and X72) xor (X41 and X62 and X73) xor (X41 and X63 and X72) xor (X42 and X61 and X72) xor (X42 and X61 and X73) xor (X42 and X62 and X71) xor (X42 and X62 and X73) xor (X42 and X63 and X71) xor (X42 and X63 and X72) xor (X43 and X61 and X72) xor (X43 and X62 and X71) xor (X43 and X62 and X73) xor (X43 and X63 and X71) xor (X43 and X63 and X73));
    F22  <= ((X02 and X12) xor (X00 and X13) xor (X02 and X13) xor (X03 and X12) xor (X22) xor (X32) xor (X12 and X32) xor (X10 and X33) xor (X12 and X33) xor (X13 and X32) xor (X10 and X20 and X33) xor (X10 and X22 and X30) xor (X10 and X22 and X32) xor (X10 and X22 and X33) xor (X10 and X23 and X30) xor (X10 and X23 and X32) xor (X12 and X20 and X32) xor (X12 and X20 and X33) xor (X12 and X23 and X30) xor (X12 and X23 and X33) xor (X13 and X20 and X30) xor (X13 and X20 and X32) xor (X13 and X20 and X33) xor (X13 and X22 and X30) xor (X13 and X22 and X32) xor (X13 and X23 and X32) xor (X42) xor (X00 and X20 and X43) xor (X00 and X22 and X40) xor (X00 and X22 and X42) xor (X00 and X22 and X43) xor (X00 and X23 and X40) xor (X00 and X23 and X42) xor (X02 and X20 and X42) xor (X02 and X20 and X43) xor (X02 and X23 and X40) xor (X02 and X23 and X43) xor (X03 and X20 and X40) xor (X03 and X20 and X42) xor (X03 and X20 and X43) xor (X03 and X22 and X40) xor (X03 and X22 and X42) xor (X03 and X23 and X42) xor (X10 and X20 and X43) xor (X10 and X22 and X40) xor (X10 and X22 and X42) xor (X10 and X22 and X43) xor (X10 and X23 and X40) xor (X10 and X23 and X42) xor (X12 and X20 and X42) xor (X12 and X20 and X43) xor (X12 and X23 and X40) xor (X12 and X23 and X43) xor (X13 and X20 and X40) xor (X13 and X20 and X42) xor (X13 and X20 and X43) xor (X13 and X22 and X40) xor (X13 and X22 and X42) xor (X13 and X23 and X42) xor (X32 and X42) xor (X30 and X43) xor (X32 and X43) xor (X33 and X42) xor (X10 and X30 and X43) xor (X10 and X32 and X40) xor (X10 and X32 and X42) xor (X10 and X32 and X43) xor (X10 and X33 and X40) xor (X10 and X33 and X42) xor (X12 and X30 and X42) xor (X12 and X30 and X43) xor (X12 and X33 and X40) xor (X12 and X33 and X43) xor (X13 and X30 and X40) xor (X13 and X30 and X42) xor (X13 and X30 and X43) xor (X13 and X32 and X40) xor (X13 and X32 and X42) xor (X13 and X33 and X42) xor (X20 and X30 and X43) xor (X20 and X32 and X40) xor (X20 and X32 and X42) xor (X20 and X32 and X43) xor (X20 and X33 and X40) xor (X20 and X33 and X42) xor (X22 and X30 and X42) xor (X22 and X30 and X43) xor (X22 and X33 and X40) xor (X22 and X33 and X43) xor (X23 and X30 and X40) xor (X23 and X30 and X42) xor (X23 and X30 and X43) xor (X23 and X32 and X40) xor (X23 and X32 and X42) xor (X23 and X33 and X42) xor (X02 and X52) xor (X00 and X53) xor (X02 and X53) xor (X03 and X52) xor (X22 and X52) xor (X20 and X53) xor (X22 and X53) xor (X23 and X52) xor (X00 and X20 and X53) xor (X00 and X22 and X50) xor (X00 and X22 and X52) xor (X00 and X22 and X53) xor (X00 and X23 and X50) xor (X00 and X23 and X52) xor (X02 and X20 and X52) xor (X02 and X20 and X53) xor (X02 and X23 and X50) xor (X02 and X23 and X53) xor (X03 and X20 and X50) xor (X03 and X20 and X52) xor (X03 and X20 and X53) xor (X03 and X22 and X50) xor (X03 and X22 and X52) xor (X03 and X23 and X52) xor (X32 and X52) xor (X30 and X53) xor (X32 and X53) xor (X33 and X52) xor (X00 and X30 and X53) xor (X00 and X32 and X50) xor (X00 and X32 and X52) xor (X00 and X32 and X53) xor (X00 and X33 and X50) xor (X00 and X33 and X52) xor (X02 and X30 and X52) xor (X02 and X30 and X53) xor (X02 and X33 and X50) xor (X02 and X33 and X53) xor (X03 and X30 and X50) xor (X03 and X30 and X52) xor (X03 and X30 and X53) xor (X03 and X32 and X50) xor (X03 and X32 and X52) xor (X03 and X33 and X52) xor (X10 and X30 and X53) xor (X10 and X32 and X50) xor (X10 and X32 and X52) xor (X10 and X32 and X53) xor (X10 and X33 and X50) xor (X10 and X33 and X52) xor (X12 and X30 and X52) xor (X12 and X30 and X53) xor (X12 and X33 and X50) xor (X12 and X33 and X53) xor (X13 and X30 and X50) xor (X13 and X30 and X52) xor (X13 and X30 and X53) xor (X13 and X32 and X50) xor (X13 and X32 and X52) xor (X13 and X33 and X52) xor (X42 and X52) xor (X40 and X53) xor (X42 and X53) xor (X43 and X52) xor (X00 and X40 and X53) xor (X00 and X42 and X50) xor (X00 and X42 and X52) xor (X00 and X42 and X53) xor (X00 and X43 and X50) xor (X00 and X43 and X52) xor (X02 and X40 and X52) xor (X02 and X40 and X53) xor (X02 and X43 and X50) xor (X02 and X43 and X53) xor (X03 and X40 and X50) xor (X03 and X40 and X52) xor (X03 and X40 and X53) xor (X03 and X42 and X50) xor (X03 and X42 and X52) xor (X03 and X43 and X52) xor (X20 and X40 and X53) xor (X20 and X42 and X50) xor (X20 and X42 and X52) xor (X20 and X42 and X53) xor (X20 and X43 and X50) xor (X20 and X43 and X52) xor (X22 and X40 and X52) xor (X22 and X40 and X53) xor (X22 and X43 and X50) xor (X22 and X43 and X53) xor (X23 and X40 and X50) xor (X23 and X40 and X52) xor (X23 and X40 and X53) xor (X23 and X42 and X50) xor (X23 and X42 and X52) xor (X23 and X43 and X52) xor (X30 and X40 and X53) xor (X30 and X42 and X50) xor (X30 and X42 and X52) xor (X30 and X42 and X53) xor (X30 and X43 and X50) xor (X30 and X43 and X52) xor (X32 and X40 and X52) xor (X32 and X40 and X53) xor (X32 and X43 and X50) xor (X32 and X43 and X53) xor (X33 and X40 and X50) xor (X33 and X40 and X52) xor (X33 and X40 and X53) xor (X33 and X42 and X50) xor (X33 and X42 and X52) xor (X33 and X43 and X52) xor (X10 and X20 and X63) xor (X10 and X22 and X60) xor (X10 and X22 and X62) xor (X10 and X22 and X63) xor (X10 and X23 and X60) xor (X10 and X23 and X62) xor (X12 and X20 and X62) xor (X12 and X20 and X63) xor (X12 and X23 and X60) xor (X12 and X23 and X63) xor (X13 and X20 and X60) xor (X13 and X20 and X62) xor (X13 and X20 and X63) xor (X13 and X22 and X60) xor (X13 and X22 and X62) xor (X13 and X23 and X62) xor (X32 and X62) xor (X30 and X63) xor (X32 and X63) xor (X33 and X62) xor (X00 and X30 and X63) xor (X00 and X32 and X60) xor (X00 and X32 and X62) xor (X00 and X32 and X63) xor (X00 and X33 and X60) xor (X00 and X33 and X62) xor (X02 and X30 and X62) xor (X02 and X30 and X63) xor (X02 and X33 and X60) xor (X02 and X33 and X63) xor (X03 and X30 and X60) xor (X03 and X30 and X62) xor (X03 and X30 and X63) xor (X03 and X32 and X60) xor (X03 and X32 and X62) xor (X03 and X33 and X62) xor (X10 and X30 and X63) xor (X10 and X32 and X60) xor (X10 and X32 and X62) xor (X10 and X32 and X63) xor (X10 and X33 and X60) xor (X10 and X33 and X62) xor (X12 and X30 and X62) xor (X12 and X30 and X63) xor (X12 and X33 and X60) xor (X12 and X33 and X63) xor (X13 and X30 and X60) xor (X13 and X30 and X62) xor (X13 and X30 and X63) xor (X13 and X32 and X60) xor (X13 and X32 and X62) xor (X13 and X33 and X62) xor (X20 and X30 and X63) xor (X20 and X32 and X60) xor (X20 and X32 and X62) xor (X20 and X32 and X63) xor (X20 and X33 and X60) xor (X20 and X33 and X62) xor (X22 and X30 and X62) xor (X22 and X30 and X63) xor (X22 and X33 and X60) xor (X22 and X33 and X63) xor (X23 and X30 and X60) xor (X23 and X30 and X62) xor (X23 and X30 and X63) xor (X23 and X32 and X60) xor (X23 and X32 and X62) xor (X23 and X33 and X62) xor (X52 and X62) xor (X50 and X63) xor (X52 and X63) xor (X53 and X62) xor (X00 and X50 and X63) xor (X00 and X52 and X60) xor (X00 and X52 and X62) xor (X00 and X52 and X63) xor (X00 and X53 and X60) xor (X00 and X53 and X62) xor (X02 and X50 and X62) xor (X02 and X50 and X63) xor (X02 and X53 and X60) xor (X02 and X53 and X63) xor (X03 and X50 and X60) xor (X03 and X50 and X62) xor (X03 and X50 and X63) xor (X03 and X52 and X60) xor (X03 and X52 and X62) xor (X03 and X53 and X62) xor (X10 and X50 and X63) xor (X10 and X52 and X60) xor (X10 and X52 and X62) xor (X10 and X52 and X63) xor (X10 and X53 and X60) xor (X10 and X53 and X62) xor (X12 and X50 and X62) xor (X12 and X50 and X63) xor (X12 and X53 and X60) xor (X12 and X53 and X63) xor (X13 and X50 and X60) xor (X13 and X50 and X62) xor (X13 and X50 and X63) xor (X13 and X52 and X60) xor (X13 and X52 and X62) xor (X13 and X53 and X62) xor (X20 and X50 and X63) xor (X20 and X52 and X60) xor (X20 and X52 and X62) xor (X20 and X52 and X63) xor (X20 and X53 and X60) xor (X20 and X53 and X62) xor (X22 and X50 and X62) xor (X22 and X50 and X63) xor (X22 and X53 and X60) xor (X22 and X53 and X63) xor (X23 and X50 and X60) xor (X23 and X50 and X62) xor (X23 and X50 and X63) xor (X23 and X52 and X60) xor (X23 and X52 and X62) xor (X23 and X53 and X62) xor (X40 and X50 and X63) xor (X40 and X52 and X60) xor (X40 and X52 and X62) xor (X40 and X52 and X63) xor (X40 and X53 and X60) xor (X40 and X53 and X62) xor (X42 and X50 and X62) xor (X42 and X50 and X63) xor (X42 and X53 and X60) xor (X42 and X53 and X63) xor (X43 and X50 and X60) xor (X43 and X50 and X62) xor (X43 and X50 and X63) xor (X43 and X52 and X60) xor (X43 and X52 and X62) xor (X43 and X53 and X62) xor (X72) xor (X12 and X72) xor (X10 and X73) xor (X12 and X73) xor (X13 and X72) xor (X00 and X10 and X73) xor (X00 and X12 and X70) xor (X00 and X12 and X72) xor (X00 and X12 and X73) xor (X00 and X13 and X70) xor (X00 and X13 and X72) xor (X02 and X10 and X72) xor (X02 and X10 and X73) xor (X02 and X13 and X70) xor (X02 and X13 and X73) xor (X03 and X10 and X70) xor (X03 and X10 and X72) xor (X03 and X10 and X73) xor (X03 and X12 and X70) xor (X03 and X12 and X72) xor (X03 and X13 and X72) xor (X10 and X20 and X73) xor (X10 and X22 and X70) xor (X10 and X22 and X72) xor (X10 and X22 and X73) xor (X10 and X23 and X70) xor (X10 and X23 and X72) xor (X12 and X20 and X72) xor (X12 and X20 and X73) xor (X12 and X23 and X70) xor (X12 and X23 and X73) xor (X13 and X20 and X70) xor (X13 and X20 and X72) xor (X13 and X20 and X73) xor (X13 and X22 and X70) xor (X13 and X22 and X72) xor (X13 and X23 and X72) xor (X32 and X72) xor (X30 and X73) xor (X32 and X73) xor (X33 and X72) xor (X00 and X30 and X73) xor (X00 and X32 and X70) xor (X00 and X32 and X72) xor (X00 and X32 and X73) xor (X00 and X33 and X70) xor (X00 and X33 and X72) xor (X02 and X30 and X72) xor (X02 and X30 and X73) xor (X02 and X33 and X70) xor (X02 and X33 and X73) xor (X03 and X30 and X70) xor (X03 and X30 and X72) xor (X03 and X30 and X73) xor (X03 and X32 and X70) xor (X03 and X32 and X72) xor (X03 and X33 and X72) xor (X42 and X72) xor (X40 and X73) xor (X42 and X73) xor (X43 and X72) xor (X00 and X40 and X73) xor (X00 and X42 and X70) xor (X00 and X42 and X72) xor (X00 and X42 and X73) xor (X00 and X43 and X70) xor (X00 and X43 and X72) xor (X02 and X40 and X72) xor (X02 and X40 and X73) xor (X02 and X43 and X70) xor (X02 and X43 and X73) xor (X03 and X40 and X70) xor (X03 and X40 and X72) xor (X03 and X40 and X73) xor (X03 and X42 and X70) xor (X03 and X42 and X72) xor (X03 and X43 and X72) xor (X10 and X40 and X73) xor (X10 and X42 and X70) xor (X10 and X42 and X72) xor (X10 and X42 and X73) xor (X10 and X43 and X70) xor (X10 and X43 and X72) xor (X12 and X40 and X72) xor (X12 and X40 and X73) xor (X12 and X43 and X70) xor (X12 and X43 and X73) xor (X13 and X40 and X70) xor (X13 and X40 and X72) xor (X13 and X40 and X73) xor (X13 and X42 and X70) xor (X13 and X42 and X72) xor (X13 and X43 and X72) xor (X30 and X40 and X73) xor (X30 and X42 and X70) xor (X30 and X42 and X72) xor (X30 and X42 and X73) xor (X30 and X43 and X70) xor (X30 and X43 and X72) xor (X32 and X40 and X72) xor (X32 and X40 and X73) xor (X32 and X43 and X70) xor (X32 and X43 and X73) xor (X33 and X40 and X70) xor (X33 and X40 and X72) xor (X33 and X40 and X73) xor (X33 and X42 and X70) xor (X33 and X42 and X72) xor (X33 and X43 and X72) xor (X52 and X72) xor (X50 and X73) xor (X52 and X73) xor (X53 and X72) xor (X00 and X50 and X73) xor (X00 and X52 and X70) xor (X00 and X52 and X72) xor (X00 and X52 and X73) xor (X00 and X53 and X70) xor (X00 and X53 and X72) xor (X02 and X50 and X72) xor (X02 and X50 and X73) xor (X02 and X53 and X70) xor (X02 and X53 and X73) xor (X03 and X50 and X70) xor (X03 and X50 and X72) xor (X03 and X50 and X73) xor (X03 and X52 and X70) xor (X03 and X52 and X72) xor (X03 and X53 and X72) xor (X10 and X50 and X73) xor (X10 and X52 and X70) xor (X10 and X52 and X72) xor (X10 and X52 and X73) xor (X10 and X53 and X70) xor (X10 and X53 and X72) xor (X12 and X50 and X72) xor (X12 and X50 and X73) xor (X12 and X53 and X70) xor (X12 and X53 and X73) xor (X13 and X50 and X70) xor (X13 and X50 and X72) xor (X13 and X50 and X73) xor (X13 and X52 and X70) xor (X13 and X52 and X72) xor (X13 and X53 and X72) xor (X62 and X72) xor (X60 and X73) xor (X62 and X73) xor (X63 and X72) xor (X00 and X60 and X73) xor (X00 and X62 and X70) xor (X00 and X62 and X72) xor (X00 and X62 and X73) xor (X00 and X63 and X70) xor (X00 and X63 and X72) xor (X02 and X60 and X72) xor (X02 and X60 and X73) xor (X02 and X63 and X70) xor (X02 and X63 and X73) xor (X03 and X60 and X70) xor (X03 and X60 and X72) xor (X03 and X60 and X73) xor (X03 and X62 and X70) xor (X03 and X62 and X72) xor (X03 and X63 and X72) xor (X10 and X60 and X73) xor (X10 and X62 and X70) xor (X10 and X62 and X72) xor (X10 and X62 and X73) xor (X10 and X63 and X70) xor (X10 and X63 and X72) xor (X12 and X60 and X72) xor (X12 and X60 and X73) xor (X12 and X63 and X70) xor (X12 and X63 and X73) xor (X13 and X60 and X70) xor (X13 and X60 and X72) xor (X13 and X60 and X73) xor (X13 and X62 and X70) xor (X13 and X62 and X72) xor (X13 and X63 and X72) xor (X40 and X60 and X73) xor (X40 and X62 and X70) xor (X40 and X62 and X72) xor (X40 and X62 and X73) xor (X40 and X63 and X70) xor (X40 and X63 and X72) xor (X42 and X60 and X72) xor (X42 and X60 and X73) xor (X42 and X63 and X70) xor (X42 and X63 and X73) xor (X43 and X60 and X70) xor (X43 and X60 and X72) xor (X43 and X60 and X73) xor (X43 and X62 and X70) xor (X43 and X62 and X72) xor (X43 and X63 and X72));
    F23  <= ((X03 and X13) xor (X03 and X10) xor (X03 and X11) xor (X0_1 and X10) xor (X23) xor (X33) xor (X13 and X33) xor (X13 and X30) xor (X13 and X31) xor (X11 and X30) xor (X10 and X20 and X31) xor (X10 and X21 and X30) xor (X10 and X21 and X33) xor (X10 and X23 and X31) xor (X10 and X23 and X33) xor (X11 and X20 and X31) xor (X11 and X20 and X33) xor (X11 and X21 and X33) xor (X11 and X23 and X30) xor (X11 and X23 and X31) xor (X11 and X23 and X33) xor (X13 and X20 and X31) xor (X13 and X21 and X30) xor (X13 and X21 and X31) xor (X13 and X21 and X33) xor (X13 and X23 and X30) xor (X43) xor (X00 and X20 and X41) xor (X00 and X21 and X40) xor (X00 and X21 and X43) xor (X00 and X23 and X41) xor (X00 and X23 and X43) xor (X0_1 and X20 and X41) xor (X0_1 and X20 and X43) xor (X0_1 and X21 and X43) xor (X0_1 and X23 and X40) xor (X0_1 and X23 and X41) xor (X0_1 and X23 and X43) xor (X03 and X20 and X41) xor (X03 and X21 and X40) xor (X03 and X21 and X41) xor (X03 and X21 and X43) xor (X03 and X23 and X40) xor (X10 and X20 and X41) xor (X10 and X21 and X40) xor (X10 and X21 and X43) xor (X10 and X23 and X41) xor (X10 and X23 and X43) xor (X11 and X20 and X41) xor (X11 and X20 and X43) xor (X11 and X21 and X43) xor (X11 and X23 and X40) xor (X11 and X23 and X41) xor (X11 and X23 and X43) xor (X13 and X20 and X41) xor (X13 and X21 and X40) xor (X13 and X21 and X41) xor (X13 and X21 and X43) xor (X13 and X23 and X40) xor (X33 and X43) xor (X33 and X40) xor (X33 and X41) xor (X31 and X40) xor (X10 and X30 and X41) xor (X10 and X31 and X40) xor (X10 and X31 and X43) xor (X10 and X33 and X41) xor (X10 and X33 and X43) xor (X11 and X30 and X41) xor (X11 and X30 and X43) xor (X11 and X31 and X43) xor (X11 and X33 and X40) xor (X11 and X33 and X41) xor (X11 and X33 and X43) xor (X13 and X30 and X41) xor (X13 and X31 and X40) xor (X13 and X31 and X41) xor (X13 and X31 and X43) xor (X13 and X33 and X40) xor (X20 and X30 and X41) xor (X20 and X31 and X40) xor (X20 and X31 and X43) xor (X20 and X33 and X41) xor (X20 and X33 and X43) xor (X21 and X30 and X41) xor (X21 and X30 and X43) xor (X21 and X31 and X43) xor (X21 and X33 and X40) xor (X21 and X33 and X41) xor (X21 and X33 and X43) xor (X23 and X30 and X41) xor (X23 and X31 and X40) xor (X23 and X31 and X41) xor (X23 and X31 and X43) xor (X23 and X33 and X40) xor (X03 and X53) xor (X03 and X50) xor (X03 and X51) xor (X0_1 and X50) xor (X23 and X53) xor (X23 and X50) xor (X23 and X51) xor (X21 and X50) xor (X00 and X20 and X51) xor (X00 and X21 and X50) xor (X00 and X21 and X53) xor (X00 and X23 and X51) xor (X00 and X23 and X53) xor (X0_1 and X20 and X51) xor (X0_1 and X20 and X53) xor (X0_1 and X21 and X53) xor (X0_1 and X23 and X50) xor (X0_1 and X23 and X51) xor (X0_1 and X23 and X53) xor (X03 and X20 and X51) xor (X03 and X21 and X50) xor (X03 and X21 and X51) xor (X03 and X21 and X53) xor (X03 and X23 and X50) xor (X33 and X53) xor (X33 and X50) xor (X33 and X51) xor (X31 and X50) xor (X00 and X30 and X51) xor (X00 and X31 and X50) xor (X00 and X31 and X53) xor (X00 and X33 and X51) xor (X00 and X33 and X53) xor (X0_1 and X30 and X51) xor (X0_1 and X30 and X53) xor (X0_1 and X31 and X53) xor (X0_1 and X33 and X50) xor (X0_1 and X33 and X51) xor (X0_1 and X33 and X53) xor (X03 and X30 and X51) xor (X03 and X31 and X50) xor (X03 and X31 and X51) xor (X03 and X31 and X53) xor (X03 and X33 and X50) xor (X10 and X30 and X51) xor (X10 and X31 and X50) xor (X10 and X31 and X53) xor (X10 and X33 and X51) xor (X10 and X33 and X53) xor (X11 and X30 and X51) xor (X11 and X30 and X53) xor (X11 and X31 and X53) xor (X11 and X33 and X50) xor (X11 and X33 and X51) xor (X11 and X33 and X53) xor (X13 and X30 and X51) xor (X13 and X31 and X50) xor (X13 and X31 and X51) xor (X13 and X31 and X53) xor (X13 and X33 and X50) xor (X43 and X53) xor (X43 and X50) xor (X43 and X51) xor (X41 and X50) xor (X00 and X40 and X51) xor (X00 and X41 and X50) xor (X00 and X41 and X53) xor (X00 and X43 and X51) xor (X00 and X43 and X53) xor (X0_1 and X40 and X51) xor (X0_1 and X40 and X53) xor (X0_1 and X41 and X53) xor (X0_1 and X43 and X50) xor (X0_1 and X43 and X51) xor (X0_1 and X43 and X53) xor (X03 and X40 and X51) xor (X03 and X41 and X50) xor (X03 and X41 and X51) xor (X03 and X41 and X53) xor (X03 and X43 and X50) xor (X20 and X40 and X51) xor (X20 and X41 and X50) xor (X20 and X41 and X53) xor (X20 and X43 and X51) xor (X20 and X43 and X53) xor (X21 and X40 and X51) xor (X21 and X40 and X53) xor (X21 and X41 and X53) xor (X21 and X43 and X50) xor (X21 and X43 and X51) xor (X21 and X43 and X53) xor (X23 and X40 and X51) xor (X23 and X41 and X50) xor (X23 and X41 and X51) xor (X23 and X41 and X53) xor (X23 and X43 and X50) xor (X30 and X40 and X51) xor (X30 and X41 and X50) xor (X30 and X41 and X53) xor (X30 and X43 and X51) xor (X30 and X43 and X53) xor (X31 and X40 and X51) xor (X31 and X40 and X53) xor (X31 and X41 and X53) xor (X31 and X43 and X50) xor (X31 and X43 and X51) xor (X31 and X43 and X53) xor (X33 and X40 and X51) xor (X33 and X41 and X50) xor (X33 and X41 and X51) xor (X33 and X41 and X53) xor (X33 and X43 and X50) xor (X10 and X20 and X61) xor (X10 and X21 and X60) xor (X10 and X21 and X63) xor (X10 and X23 and X61) xor (X10 and X23 and X63) xor (X11 and X20 and X61) xor (X11 and X20 and X63) xor (X11 and X21 and X63) xor (X11 and X23 and X60) xor (X11 and X23 and X61) xor (X11 and X23 and X63) xor (X13 and X20 and X61) xor (X13 and X21 and X60) xor (X13 and X21 and X61) xor (X13 and X21 and X63) xor (X13 and X23 and X60) xor (X33 and X63) xor (X33 and X60) xor (X33 and X61) xor (X31 and X60) xor (X00 and X30 and X61) xor (X00 and X31 and X60) xor (X00 and X31 and X63) xor (X00 and X33 and X61) xor (X00 and X33 and X63) xor (X0_1 and X30 and X61) xor (X0_1 and X30 and X63) xor (X0_1 and X31 and X63) xor (X0_1 and X33 and X60) xor (X0_1 and X33 and X61) xor (X0_1 and X33 and X63) xor (X03 and X30 and X61) xor (X03 and X31 and X60) xor (X03 and X31 and X61) xor (X03 and X31 and X63) xor (X03 and X33 and X60) xor (X10 and X30 and X61) xor (X10 and X31 and X60) xor (X10 and X31 and X63) xor (X10 and X33 and X61) xor (X10 and X33 and X63) xor (X11 and X30 and X61) xor (X11 and X30 and X63) xor (X11 and X31 and X63) xor (X11 and X33 and X60) xor (X11 and X33 and X61) xor (X11 and X33 and X63) xor (X13 and X30 and X61) xor (X13 and X31 and X60) xor (X13 and X31 and X61) xor (X13 and X31 and X63) xor (X13 and X33 and X60) xor (X20 and X30 and X61) xor (X20 and X31 and X60) xor (X20 and X31 and X63) xor (X20 and X33 and X61) xor (X20 and X33 and X63) xor (X21 and X30 and X61) xor (X21 and X30 and X63) xor (X21 and X31 and X63) xor (X21 and X33 and X60) xor (X21 and X33 and X61) xor (X21 and X33 and X63) xor (X23 and X30 and X61) xor (X23 and X31 and X60) xor (X23 and X31 and X61) xor (X23 and X31 and X63) xor (X23 and X33 and X60) xor (X53 and X63) xor (X53 and X60) xor (X53 and X61) xor (X51 and X60) xor (X00 and X50 and X61) xor (X00 and X51 and X60) xor (X00 and X51 and X63) xor (X00 and X53 and X61) xor (X00 and X53 and X63) xor (X0_1 and X50 and X61) xor (X0_1 and X50 and X63) xor (X0_1 and X51 and X63) xor (X0_1 and X53 and X60) xor (X0_1 and X53 and X61) xor (X0_1 and X53 and X63) xor (X03 and X50 and X61) xor (X03 and X51 and X60) xor (X03 and X51 and X61) xor (X03 and X51 and X63) xor (X03 and X53 and X60) xor (X10 and X50 and X61) xor (X10 and X51 and X60) xor (X10 and X51 and X63) xor (X10 and X53 and X61) xor (X10 and X53 and X63) xor (X11 and X50 and X61) xor (X11 and X50 and X63) xor (X11 and X51 and X63) xor (X11 and X53 and X60) xor (X11 and X53 and X61) xor (X11 and X53 and X63) xor (X13 and X50 and X61) xor (X13 and X51 and X60) xor (X13 and X51 and X61) xor (X13 and X51 and X63) xor (X13 and X53 and X60) xor (X20 and X50 and X61) xor (X20 and X51 and X60) xor (X20 and X51 and X63) xor (X20 and X53 and X61) xor (X20 and X53 and X63) xor (X21 and X50 and X61) xor (X21 and X50 and X63) xor (X21 and X51 and X63) xor (X21 and X53 and X60) xor (X21 and X53 and X61) xor (X21 and X53 and X63) xor (X23 and X50 and X61) xor (X23 and X51 and X60) xor (X23 and X51 and X61) xor (X23 and X51 and X63) xor (X23 and X53 and X60) xor (X40 and X50 and X61) xor (X40 and X51 and X60) xor (X40 and X51 and X63) xor (X40 and X53 and X61) xor (X40 and X53 and X63) xor (X41 and X50 and X61) xor (X41 and X50 and X63) xor (X41 and X51 and X63) xor (X41 and X53 and X60) xor (X41 and X53 and X61) xor (X41 and X53 and X63) xor (X43 and X50 and X61) xor (X43 and X51 and X60) xor (X43 and X51 and X61) xor (X43 and X51 and X63) xor (X43 and X53 and X60) xor (X73) xor (X13 and X73) xor (X13 and X70) xor (X13 and X71) xor (X11 and X70) xor (X00 and X10 and X71) xor (X00 and X11 and X70) xor (X00 and X11 and X73) xor (X00 and X13 and X71) xor (X00 and X13 and X73) xor (X0_1 and X10 and X71) xor (X0_1 and X10 and X73) xor (X0_1 and X11 and X73) xor (X0_1 and X13 and X70) xor (X0_1 and X13 and X71) xor (X0_1 and X13 and X73) xor (X03 and X10 and X71) xor (X03 and X11 and X70) xor (X03 and X11 and X71) xor (X03 and X11 and X73) xor (X03 and X13 and X70) xor (X10 and X20 and X71) xor (X10 and X21 and X70) xor (X10 and X21 and X73) xor (X10 and X23 and X71) xor (X10 and X23 and X73) xor (X11 and X20 and X71) xor (X11 and X20 and X73) xor (X11 and X21 and X73) xor (X11 and X23 and X70) xor (X11 and X23 and X71) xor (X11 and X23 and X73) xor (X13 and X20 and X71) xor (X13 and X21 and X70) xor (X13 and X21 and X71) xor (X13 and X21 and X73) xor (X13 and X23 and X70) xor (X33 and X73) xor (X33 and X70) xor (X33 and X71) xor (X31 and X70) xor (X00 and X30 and X71) xor (X00 and X31 and X70) xor (X00 and X31 and X73) xor (X00 and X33 and X71) xor (X00 and X33 and X73) xor (X0_1 and X30 and X71) xor (X0_1 and X30 and X73) xor (X0_1 and X31 and X73) xor (X0_1 and X33 and X70) xor (X0_1 and X33 and X71) xor (X0_1 and X33 and X73) xor (X03 and X30 and X71) xor (X03 and X31 and X70) xor (X03 and X31 and X71) xor (X03 and X31 and X73) xor (X03 and X33 and X70) xor (X43 and X73) xor (X43 and X70) xor (X43 and X71) xor (X41 and X70) xor (X00 and X40 and X71) xor (X00 and X41 and X70) xor (X00 and X41 and X73) xor (X00 and X43 and X71) xor (X00 and X43 and X73) xor (X0_1 and X40 and X71) xor (X0_1 and X40 and X73) xor (X0_1 and X41 and X73) xor (X0_1 and X43 and X70) xor (X0_1 and X43 and X71) xor (X0_1 and X43 and X73) xor (X03 and X40 and X71) xor (X03 and X41 and X70) xor (X03 and X41 and X71) xor (X03 and X41 and X73) xor (X03 and X43 and X70) xor (X10 and X40 and X71) xor (X10 and X41 and X70) xor (X10 and X41 and X73) xor (X10 and X43 and X71) xor (X10 and X43 and X73) xor (X11 and X40 and X71) xor (X11 and X40 and X73) xor (X11 and X41 and X73) xor (X11 and X43 and X70) xor (X11 and X43 and X71) xor (X11 and X43 and X73) xor (X13 and X40 and X71) xor (X13 and X41 and X70) xor (X13 and X41 and X71) xor (X13 and X41 and X73) xor (X13 and X43 and X70) xor (X30 and X40 and X71) xor (X30 and X41 and X70) xor (X30 and X41 and X73) xor (X30 and X43 and X71) xor (X30 and X43 and X73) xor (X31 and X40 and X71) xor (X31 and X40 and X73) xor (X31 and X41 and X73) xor (X31 and X43 and X70) xor (X31 and X43 and X71) xor (X31 and X43 and X73) xor (X33 and X40 and X71) xor (X33 and X41 and X70) xor (X33 and X41 and X71) xor (X33 and X41 and X73) xor (X33 and X43 and X70) xor (X53 and X73) xor (X53 and X70) xor (X53 and X71) xor (X51 and X70) xor (X00 and X50 and X71) xor (X00 and X51 and X70) xor (X00 and X51 and X73) xor (X00 and X53 and X71) xor (X00 and X53 and X73) xor (X0_1 and X50 and X71) xor (X0_1 and X50 and X73) xor (X0_1 and X51 and X73) xor (X0_1 and X53 and X70) xor (X0_1 and X53 and X71) xor (X0_1 and X53 and X73) xor (X03 and X50 and X71) xor (X03 and X51 and X70) xor (X03 and X51 and X71) xor (X03 and X51 and X73) xor (X03 and X53 and X70) xor (X10 and X50 and X71) xor (X10 and X51 and X70) xor (X10 and X51 and X73) xor (X10 and X53 and X71) xor (X10 and X53 and X73) xor (X11 and X50 and X71) xor (X11 and X50 and X73) xor (X11 and X51 and X73) xor (X11 and X53 and X70) xor (X11 and X53 and X71) xor (X11 and X53 and X73) xor (X13 and X50 and X71) xor (X13 and X51 and X70) xor (X13 and X51 and X71) xor (X13 and X51 and X73) xor (X13 and X53 and X70) xor (X63 and X73) xor (X63 and X70) xor (X63 and X71) xor (X61 and X70) xor (X00 and X60 and X71) xor (X00 and X61 and X70) xor (X00 and X61 and X73) xor (X00 and X63 and X71) xor (X00 and X63 and X73) xor (X0_1 and X60 and X71) xor (X0_1 and X60 and X73) xor (X0_1 and X61 and X73) xor (X0_1 and X63 and X70) xor (X0_1 and X63 and X71) xor (X0_1 and X63 and X73) xor (X03 and X60 and X71) xor (X03 and X61 and X70) xor (X03 and X61 and X71) xor (X03 and X61 and X73) xor (X03 and X63 and X70) xor (X10 and X60 and X71) xor (X10 and X61 and X70) xor (X10 and X61 and X73) xor (X10 and X63 and X71) xor (X10 and X63 and X73) xor (X11 and X60 and X71) xor (X11 and X60 and X73) xor (X11 and X61 and X73) xor (X11 and X63 and X70) xor (X11 and X63 and X71) xor (X11 and X63 and X73) xor (X13 and X60 and X71) xor (X13 and X61 and X70) xor (X13 and X61 and X71) xor (X13 and X61 and X73) xor (X13 and X63 and X70) xor (X40 and X60 and X71) xor (X40 and X61 and X70) xor (X40 and X61 and X73) xor (X40 and X63 and X71) xor (X40 and X63 and X73) xor (X41 and X60 and X71) xor (X41 and X60 and X73) xor (X41 and X61 and X73) xor (X41 and X63 and X70) xor (X41 and X63 and X71) xor (X41 and X63 and X73) xor (X43 and X60 and X71) xor (X43 and X61 and X70) xor (X43 and X61 and X71) xor (X43 and X61 and X73) xor (X43 and X63 and X70));
    F30  <= ((X10) xor (X00 and X10) xor (X00 and X11) xor (X02 and X10) xor (X00 and X12) xor (X10 and X20) xor (X10 and X21) xor (X12 and X20) xor (X10 and X22) xor (X00 and X10 and X20) xor (X00 and X10 and X22) xor (X00 and X11 and X21) xor (X00 and X11 and X22) xor (X00 and X12 and X21) xor (X0_1 and X10 and X20) xor (X0_1 and X10 and X22) xor (X0_1 and X11 and X20) xor (X0_1 and X12 and X20) xor (X0_1 and X12 and X21) xor (X02 and X10 and X20) xor (X02 and X10 and X21) xor (X02 and X11 and X20) xor (X02 and X11 and X21) xor (X02 and X12 and X20) xor (X02 and X12 and X22) xor (X30) xor (X00 and X10 and X30) xor (X00 and X10 and X32) xor (X00 and X11 and X31) xor (X00 and X11 and X32) xor (X00 and X12 and X31) xor (X0_1 and X10 and X30) xor (X0_1 and X10 and X32) xor (X0_1 and X11 and X30) xor (X0_1 and X12 and X30) xor (X0_1 and X12 and X31) xor (X02 and X10 and X30) xor (X02 and X10 and X31) xor (X02 and X11 and X30) xor (X02 and X11 and X31) xor (X02 and X12 and X30) xor (X02 and X12 and X32) xor (X20 and X30) xor (X20 and X31) xor (X22 and X30) xor (X20 and X32) xor (X40) xor (X00 and X40) xor (X00 and X41) xor (X02 and X40) xor (X00 and X42) xor (X00 and X10 and X40) xor (X00 and X10 and X42) xor (X00 and X11 and X41) xor (X00 and X11 and X42) xor (X00 and X12 and X41) xor (X0_1 and X10 and X40) xor (X0_1 and X10 and X42) xor (X0_1 and X11 and X40) xor (X0_1 and X12 and X40) xor (X0_1 and X12 and X41) xor (X02 and X10 and X40) xor (X02 and X10 and X41) xor (X02 and X11 and X40) xor (X02 and X11 and X41) xor (X02 and X12 and X40) xor (X02 and X12 and X42) xor (X20 and X40) xor (X20 and X41) xor (X22 and X40) xor (X20 and X42) xor (X00 and X20 and X40) xor (X00 and X20 and X42) xor (X00 and X21 and X41) xor (X00 and X21 and X42) xor (X00 and X22 and X41) xor (X0_1 and X20 and X40) xor (X0_1 and X20 and X42) xor (X0_1 and X21 and X40) xor (X0_1 and X22 and X40) xor (X0_1 and X22 and X41) xor (X02 and X20 and X40) xor (X02 and X20 and X41) xor (X02 and X21 and X40) xor (X02 and X21 and X41) xor (X02 and X22 and X40) xor (X02 and X22 and X42) xor (X10 and X20 and X40) xor (X10 and X20 and X42) xor (X10 and X21 and X41) xor (X10 and X21 and X42) xor (X10 and X22 and X41) xor (X11 and X20 and X40) xor (X11 and X20 and X42) xor (X11 and X21 and X40) xor (X11 and X22 and X40) xor (X11 and X22 and X41) xor (X12 and X20 and X40) xor (X12 and X20 and X41) xor (X12 and X21 and X40) xor (X12 and X21 and X41) xor (X12 and X22 and X40) xor (X12 and X22 and X42) xor (X30 and X40) xor (X30 and X41) xor (X32 and X40) xor (X30 and X42) xor (X10 and X50) xor (X10 and X51) xor (X12 and X50) xor (X10 and X52) xor (X20 and X50) xor (X20 and X51) xor (X22 and X50) xor (X20 and X52) xor (X20 and X30 and X50) xor (X20 and X30 and X52) xor (X20 and X31 and X51) xor (X20 and X31 and X52) xor (X20 and X32 and X51) xor (X21 and X30 and X50) xor (X21 and X30 and X52) xor (X21 and X31 and X50) xor (X21 and X32 and X50) xor (X21 and X32 and X51) xor (X22 and X30 and X50) xor (X22 and X30 and X51) xor (X22 and X31 and X50) xor (X22 and X31 and X51) xor (X22 and X32 and X50) xor (X22 and X32 and X52) xor (X00 and X40 and X50) xor (X00 and X40 and X52) xor (X00 and X41 and X51) xor (X00 and X41 and X52) xor (X00 and X42 and X51) xor (X0_1 and X40 and X50) xor (X0_1 and X40 and X52) xor (X0_1 and X41 and X50) xor (X0_1 and X42 and X50) xor (X0_1 and X42 and X51) xor (X02 and X40 and X50) xor (X02 and X40 and X51) xor (X02 and X41 and X50) xor (X02 and X41 and X51) xor (X02 and X42 and X50) xor (X02 and X42 and X52) xor (X10 and X40 and X50) xor (X10 and X40 and X52) xor (X10 and X41 and X51) xor (X10 and X41 and X52) xor (X10 and X42 and X51) xor (X11 and X40 and X50) xor (X11 and X40 and X52) xor (X11 and X41 and X50) xor (X11 and X42 and X50) xor (X11 and X42 and X51) xor (X12 and X40 and X50) xor (X12 and X40 and X51) xor (X12 and X41 and X50) xor (X12 and X41 and X51) xor (X12 and X42 and X50) xor (X12 and X42 and X52) xor (X30 and X40 and X50) xor (X30 and X40 and X52) xor (X30 and X41 and X51) xor (X30 and X41 and X52) xor (X30 and X42 and X51) xor (X31 and X40 and X50) xor (X31 and X40 and X52) xor (X31 and X41 and X50) xor (X31 and X42 and X50) xor (X31 and X42 and X51) xor (X32 and X40 and X50) xor (X32 and X40 and X51) xor (X32 and X41 and X50) xor (X32 and X41 and X51) xor (X32 and X42 and X50) xor (X32 and X42 and X52) xor (X60) xor (X00 and X60) xor (X00 and X61) xor (X02 and X60) xor (X00 and X62) xor (X00 and X10 and X60) xor (X00 and X10 and X62) xor (X00 and X11 and X61) xor (X00 and X11 and X62) xor (X00 and X12 and X61) xor (X0_1 and X10 and X60) xor (X0_1 and X10 and X62) xor (X0_1 and X11 and X60) xor (X0_1 and X12 and X60) xor (X0_1 and X12 and X61) xor (X02 and X10 and X60) xor (X02 and X10 and X61) xor (X02 and X11 and X60) xor (X02 and X11 and X61) xor (X02 and X12 and X60) xor (X02 and X12 and X62) xor (X20 and X60) xor (X20 and X61) xor (X22 and X60) xor (X20 and X62) xor (X10 and X20 and X60) xor (X10 and X20 and X62) xor (X10 and X21 and X61) xor (X10 and X21 and X62) xor (X10 and X22 and X61) xor (X11 and X20 and X60) xor (X11 and X20 and X62) xor (X11 and X21 and X60) xor (X11 and X22 and X60) xor (X11 and X22 and X61) xor (X12 and X20 and X60) xor (X12 and X20 and X61) xor (X12 and X21 and X60) xor (X12 and X21 and X61) xor (X12 and X22 and X60) xor (X12 and X22 and X62) xor (X30 and X60) xor (X30 and X61) xor (X32 and X60) xor (X30 and X62) xor (X00 and X30 and X60) xor (X00 and X30 and X62) xor (X00 and X31 and X61) xor (X00 and X31 and X62) xor (X00 and X32 and X61) xor (X0_1 and X30 and X60) xor (X0_1 and X30 and X62) xor (X0_1 and X31 and X60) xor (X0_1 and X32 and X60) xor (X0_1 and X32 and X61) xor (X02 and X30 and X60) xor (X02 and X30 and X61) xor (X02 and X31 and X60) xor (X02 and X31 and X61) xor (X02 and X32 and X60) xor (X02 and X32 and X62) xor (X40 and X60) xor (X40 and X61) xor (X42 and X60) xor (X40 and X62) xor (X10 and X40 and X60) xor (X10 and X40 and X62) xor (X10 and X41 and X61) xor (X10 and X41 and X62) xor (X10 and X42 and X61) xor (X11 and X40 and X60) xor (X11 and X40 and X62) xor (X11 and X41 and X60) xor (X11 and X42 and X60) xor (X11 and X42 and X61) xor (X12 and X40 and X60) xor (X12 and X40 and X61) xor (X12 and X41 and X60) xor (X12 and X41 and X61) xor (X12 and X42 and X60) xor (X12 and X42 and X62) xor (X50 and X60) xor (X50 and X61) xor (X52 and X60) xor (X50 and X62) xor (X00 and X50 and X60) xor (X00 and X50 and X62) xor (X00 and X51 and X61) xor (X00 and X51 and X62) xor (X00 and X52 and X61) xor (X0_1 and X50 and X60) xor (X0_1 and X50 and X62) xor (X0_1 and X51 and X60) xor (X0_1 and X52 and X60) xor (X0_1 and X52 and X61) xor (X02 and X50 and X60) xor (X02 and X50 and X61) xor (X02 and X51 and X60) xor (X02 and X51 and X61) xor (X02 and X52 and X60) xor (X02 and X52 and X62) xor (X10 and X50 and X60) xor (X10 and X50 and X62) xor (X10 and X51 and X61) xor (X10 and X51 and X62) xor (X10 and X52 and X61) xor (X11 and X50 and X60) xor (X11 and X50 and X62) xor (X11 and X51 and X60) xor (X11 and X52 and X60) xor (X11 and X52 and X61) xor (X12 and X50 and X60) xor (X12 and X50 and X61) xor (X12 and X51 and X60) xor (X12 and X51 and X61) xor (X12 and X52 and X60) xor (X12 and X52 and X62) xor (X20 and X50 and X60) xor (X20 and X50 and X62) xor (X20 and X51 and X61) xor (X20 and X51 and X62) xor (X20 and X52 and X61) xor (X21 and X50 and X60) xor (X21 and X50 and X62) xor (X21 and X51 and X60) xor (X21 and X52 and X60) xor (X21 and X52 and X61) xor (X22 and X50 and X60) xor (X22 and X50 and X61) xor (X22 and X51 and X60) xor (X22 and X51 and X61) xor (X22 and X52 and X60) xor (X22 and X52 and X62) xor (X30 and X50 and X60) xor (X30 and X50 and X62) xor (X30 and X51 and X61) xor (X30 and X51 and X62) xor (X30 and X52 and X61) xor (X31 and X50 and X60) xor (X31 and X50 and X62) xor (X31 and X51 and X60) xor (X31 and X52 and X60) xor (X31 and X52 and X61) xor (X32 and X50 and X60) xor (X32 and X50 and X61) xor (X32 and X51 and X60) xor (X32 and X51 and X61) xor (X32 and X52 and X60) xor (X32 and X52 and X62) xor (X40 and X50 and X60) xor (X40 and X50 and X62) xor (X40 and X51 and X61) xor (X40 and X51 and X62) xor (X40 and X52 and X61) xor (X41 and X50 and X60) xor (X41 and X50 and X62) xor (X41 and X51 and X60) xor (X41 and X52 and X60) xor (X41 and X52 and X61) xor (X42 and X50 and X60) xor (X42 and X50 and X61) xor (X42 and X51 and X60) xor (X42 and X51 and X61) xor (X42 and X52 and X60) xor (X42 and X52 and X62) xor (X70) xor (X00 and X20 and X70) xor (X00 and X20 and X72) xor (X00 and X21 and X71) xor (X00 and X21 and X72) xor (X00 and X22 and X71) xor (X0_1 and X20 and X70) xor (X0_1 and X20 and X72) xor (X0_1 and X21 and X70) xor (X0_1 and X22 and X70) xor (X0_1 and X22 and X71) xor (X02 and X20 and X70) xor (X02 and X20 and X71) xor (X02 and X21 and X70) xor (X02 and X21 and X71) xor (X02 and X22 and X70) xor (X02 and X22 and X72) xor (X10 and X30 and X70) xor (X10 and X30 and X72) xor (X10 and X31 and X71) xor (X10 and X31 and X72) xor (X10 and X32 and X71) xor (X11 and X30 and X70) xor (X11 and X30 and X72) xor (X11 and X31 and X70) xor (X11 and X32 and X70) xor (X11 and X32 and X71) xor (X12 and X30 and X70) xor (X12 and X30 and X71) xor (X12 and X31 and X70) xor (X12 and X31 and X71) xor (X12 and X32 and X70) xor (X12 and X32 and X72) xor (X00 and X40 and X70) xor (X00 and X40 and X72) xor (X00 and X41 and X71) xor (X00 and X41 and X72) xor (X00 and X42 and X71) xor (X0_1 and X40 and X70) xor (X0_1 and X40 and X72) xor (X0_1 and X41 and X70) xor (X0_1 and X42 and X70) xor (X0_1 and X42 and X71) xor (X02 and X40 and X70) xor (X02 and X40 and X71) xor (X02 and X41 and X70) xor (X02 and X41 and X71) xor (X02 and X42 and X70) xor (X02 and X42 and X72) xor (X50 and X70) xor (X50 and X71) xor (X52 and X70) xor (X50 and X72) xor (X00 and X50 and X70) xor (X00 and X50 and X72) xor (X00 and X51 and X71) xor (X00 and X51 and X72) xor (X00 and X52 and X71) xor (X0_1 and X50 and X70) xor (X0_1 and X50 and X72) xor (X0_1 and X51 and X70) xor (X0_1 and X52 and X70) xor (X0_1 and X52 and X71) xor (X02 and X50 and X70) xor (X02 and X50 and X71) xor (X02 and X51 and X70) xor (X02 and X51 and X71) xor (X02 and X52 and X70) xor (X02 and X52 and X72) xor (X10 and X50 and X70) xor (X10 and X50 and X72) xor (X10 and X51 and X71) xor (X10 and X51 and X72) xor (X10 and X52 and X71) xor (X11 and X50 and X70) xor (X11 and X50 and X72) xor (X11 and X51 and X70) xor (X11 and X52 and X70) xor (X11 and X52 and X71) xor (X12 and X50 and X70) xor (X12 and X50 and X71) xor (X12 and X51 and X70) xor (X12 and X51 and X71) xor (X12 and X52 and X70) xor (X12 and X52 and X72) xor (X30 and X50 and X70) xor (X30 and X50 and X72) xor (X30 and X51 and X71) xor (X30 and X51 and X72) xor (X30 and X52 and X71) xor (X31 and X50 and X70) xor (X31 and X50 and X72) xor (X31 and X51 and X70) xor (X31 and X52 and X70) xor (X31 and X52 and X71) xor (X32 and X50 and X70) xor (X32 and X50 and X71) xor (X32 and X51 and X70) xor (X32 and X51 and X71) xor (X32 and X52 and X70) xor (X32 and X52 and X72) xor (X00 and X60 and X70) xor (X00 and X60 and X72) xor (X00 and X61 and X71) xor (X00 and X61 and X72) xor (X00 and X62 and X71) xor (X0_1 and X60 and X70) xor (X0_1 and X60 and X72) xor (X0_1 and X61 and X70) xor (X0_1 and X62 and X70) xor (X0_1 and X62 and X71) xor (X02 and X60 and X70) xor (X02 and X60 and X71) xor (X02 and X61 and X70) xor (X02 and X61 and X71) xor (X02 and X62 and X70) xor (X02 and X62 and X72) xor (X20 and X60 and X70) xor (X20 and X60 and X72) xor (X20 and X61 and X71) xor (X20 and X61 and X72) xor (X20 and X62 and X71) xor (X21 and X60 and X70) xor (X21 and X60 and X72) xor (X21 and X61 and X70) xor (X21 and X62 and X70) xor (X21 and X62 and X71) xor (X22 and X60 and X70) xor (X22 and X60 and X71) xor (X22 and X61 and X70) xor (X22 and X61 and X71) xor (X22 and X62 and X70) xor (X22 and X62 and X72) xor (X40 and X60 and X70) xor (X40 and X60 and X72) xor (X40 and X61 and X71) xor (X40 and X61 and X72) xor (X40 and X62 and X71) xor (X41 and X60 and X70) xor (X41 and X60 and X72) xor (X41 and X61 and X70) xor (X41 and X62 and X70) xor (X41 and X62 and X71) xor (X42 and X60 and X70) xor (X42 and X60 and X71) xor (X42 and X61 and X70) xor (X42 and X61 and X71) xor (X42 and X62 and X70) xor (X42 and X62 and X72));
    F31  <= ((X11) xor (X0_1 and X11) xor (X0_1 and X12) xor (X02 and X11) xor (X0_1 and X13) xor (X11 and X21) xor (X11 and X22) xor (X12 and X21) xor (X11 and X23) xor (X0_1 and X11 and X21) xor (X0_1 and X11 and X22) xor (X0_1 and X12 and X22) xor (X0_1 and X12 and X23) xor (X0_1 and X13 and X22) xor (X02 and X11 and X22) xor (X02 and X11 and X23) xor (X02 and X12 and X21) xor (X02 and X12 and X23) xor (X02 and X13 and X21) xor (X02 and X13 and X22) xor (X03 and X11 and X22) xor (X03 and X12 and X21) xor (X03 and X12 and X23) xor (X03 and X13 and X21) xor (X03 and X13 and X23) xor (X31) xor (X0_1 and X11 and X31) xor (X0_1 and X11 and X32) xor (X0_1 and X12 and X32) xor (X0_1 and X12 and X33) xor (X0_1 and X13 and X32) xor (X02 and X11 and X32) xor (X02 and X11 and X33) xor (X02 and X12 and X31) xor (X02 and X12 and X33) xor (X02 and X13 and X31) xor (X02 and X13 and X32) xor (X03 and X11 and X32) xor (X03 and X12 and X31) xor (X03 and X12 and X33) xor (X03 and X13 and X31) xor (X03 and X13 and X33) xor (X21 and X31) xor (X21 and X32) xor (X22 and X31) xor (X21 and X33) xor (X41) xor (X0_1 and X41) xor (X0_1 and X42) xor (X02 and X41) xor (X0_1 and X43) xor (X0_1 and X11 and X41) xor (X0_1 and X11 and X42) xor (X0_1 and X12 and X42) xor (X0_1 and X12 and X43) xor (X0_1 and X13 and X42) xor (X02 and X11 and X42) xor (X02 and X11 and X43) xor (X02 and X12 and X41) xor (X02 and X12 and X43) xor (X02 and X13 and X41) xor (X02 and X13 and X42) xor (X03 and X11 and X42) xor (X03 and X12 and X41) xor (X03 and X12 and X43) xor (X03 and X13 and X41) xor (X03 and X13 and X43) xor (X21 and X41) xor (X21 and X42) xor (X22 and X41) xor (X21 and X43) xor (X0_1 and X21 and X41) xor (X0_1 and X21 and X42) xor (X0_1 and X22 and X42) xor (X0_1 and X22 and X43) xor (X0_1 and X23 and X42) xor (X02 and X21 and X42) xor (X02 and X21 and X43) xor (X02 and X22 and X41) xor (X02 and X22 and X43) xor (X02 and X23 and X41) xor (X02 and X23 and X42) xor (X03 and X21 and X42) xor (X03 and X22 and X41) xor (X03 and X22 and X43) xor (X03 and X23 and X41) xor (X03 and X23 and X43) xor (X11 and X21 and X41) xor (X11 and X21 and X42) xor (X11 and X22 and X42) xor (X11 and X22 and X43) xor (X11 and X23 and X42) xor (X12 and X21 and X42) xor (X12 and X21 and X43) xor (X12 and X22 and X41) xor (X12 and X22 and X43) xor (X12 and X23 and X41) xor (X12 and X23 and X42) xor (X13 and X21 and X42) xor (X13 and X22 and X41) xor (X13 and X22 and X43) xor (X13 and X23 and X41) xor (X13 and X23 and X43) xor (X31 and X41) xor (X31 and X42) xor (X32 and X41) xor (X31 and X43) xor (X11 and X51) xor (X11 and X52) xor (X12 and X51) xor (X11 and X53) xor (X21 and X51) xor (X21 and X52) xor (X22 and X51) xor (X21 and X53) xor (X21 and X31 and X51) xor (X21 and X31 and X52) xor (X21 and X32 and X52) xor (X21 and X32 and X53) xor (X21 and X33 and X52) xor (X22 and X31 and X52) xor (X22 and X31 and X53) xor (X22 and X32 and X51) xor (X22 and X32 and X53) xor (X22 and X33 and X51) xor (X22 and X33 and X52) xor (X23 and X31 and X52) xor (X23 and X32 and X51) xor (X23 and X32 and X53) xor (X23 and X33 and X51) xor (X23 and X33 and X53) xor (X0_1 and X41 and X51) xor (X0_1 and X41 and X52) xor (X0_1 and X42 and X52) xor (X0_1 and X42 and X53) xor (X0_1 and X43 and X52) xor (X02 and X41 and X52) xor (X02 and X41 and X53) xor (X02 and X42 and X51) xor (X02 and X42 and X53) xor (X02 and X43 and X51) xor (X02 and X43 and X52) xor (X03 and X41 and X52) xor (X03 and X42 and X51) xor (X03 and X42 and X53) xor (X03 and X43 and X51) xor (X03 and X43 and X53) xor (X11 and X41 and X51) xor (X11 and X41 and X52) xor (X11 and X42 and X52) xor (X11 and X42 and X53) xor (X11 and X43 and X52) xor (X12 and X41 and X52) xor (X12 and X41 and X53) xor (X12 and X42 and X51) xor (X12 and X42 and X53) xor (X12 and X43 and X51) xor (X12 and X43 and X52) xor (X13 and X41 and X52) xor (X13 and X42 and X51) xor (X13 and X42 and X53) xor (X13 and X43 and X51) xor (X13 and X43 and X53) xor (X31 and X41 and X51) xor (X31 and X41 and X52) xor (X31 and X42 and X52) xor (X31 and X42 and X53) xor (X31 and X43 and X52) xor (X32 and X41 and X52) xor (X32 and X41 and X53) xor (X32 and X42 and X51) xor (X32 and X42 and X53) xor (X32 and X43 and X51) xor (X32 and X43 and X52) xor (X33 and X41 and X52) xor (X33 and X42 and X51) xor (X33 and X42 and X53) xor (X33 and X43 and X51) xor (X33 and X43 and X53) xor (X61) xor (X0_1 and X61) xor (X0_1 and X62) xor (X02 and X61) xor (X0_1 and X63) xor (X0_1 and X11 and X61) xor (X0_1 and X11 and X62) xor (X0_1 and X12 and X62) xor (X0_1 and X12 and X63) xor (X0_1 and X13 and X62) xor (X02 and X11 and X62) xor (X02 and X11 and X63) xor (X02 and X12 and X61) xor (X02 and X12 and X63) xor (X02 and X13 and X61) xor (X02 and X13 and X62) xor (X03 and X11 and X62) xor (X03 and X12 and X61) xor (X03 and X12 and X63) xor (X03 and X13 and X61) xor (X03 and X13 and X63) xor (X21 and X61) xor (X21 and X62) xor (X22 and X61) xor (X21 and X63) xor (X11 and X21 and X61) xor (X11 and X21 and X62) xor (X11 and X22 and X62) xor (X11 and X22 and X63) xor (X11 and X23 and X62) xor (X12 and X21 and X62) xor (X12 and X21 and X63) xor (X12 and X22 and X61) xor (X12 and X22 and X63) xor (X12 and X23 and X61) xor (X12 and X23 and X62) xor (X13 and X21 and X62) xor (X13 and X22 and X61) xor (X13 and X22 and X63) xor (X13 and X23 and X61) xor (X13 and X23 and X63) xor (X31 and X61) xor (X31 and X62) xor (X32 and X61) xor (X31 and X63) xor (X0_1 and X31 and X61) xor (X0_1 and X31 and X62) xor (X0_1 and X32 and X62) xor (X0_1 and X32 and X63) xor (X0_1 and X33 and X62) xor (X02 and X31 and X62) xor (X02 and X31 and X63) xor (X02 and X32 and X61) xor (X02 and X32 and X63) xor (X02 and X33 and X61) xor (X02 and X33 and X62) xor (X03 and X31 and X62) xor (X03 and X32 and X61) xor (X03 and X32 and X63) xor (X03 and X33 and X61) xor (X03 and X33 and X63) xor (X41 and X61) xor (X41 and X62) xor (X42 and X61) xor (X41 and X63) xor (X11 and X41 and X61) xor (X11 and X41 and X62) xor (X11 and X42 and X62) xor (X11 and X42 and X63) xor (X11 and X43 and X62) xor (X12 and X41 and X62) xor (X12 and X41 and X63) xor (X12 and X42 and X61) xor (X12 and X42 and X63) xor (X12 and X43 and X61) xor (X12 and X43 and X62) xor (X13 and X41 and X62) xor (X13 and X42 and X61) xor (X13 and X42 and X63) xor (X13 and X43 and X61) xor (X13 and X43 and X63) xor (X51 and X61) xor (X51 and X62) xor (X52 and X61) xor (X51 and X63) xor (X0_1 and X51 and X61) xor (X0_1 and X51 and X62) xor (X0_1 and X52 and X62) xor (X0_1 and X52 and X63) xor (X0_1 and X53 and X62) xor (X02 and X51 and X62) xor (X02 and X51 and X63) xor (X02 and X52 and X61) xor (X02 and X52 and X63) xor (X02 and X53 and X61) xor (X02 and X53 and X62) xor (X03 and X51 and X62) xor (X03 and X52 and X61) xor (X03 and X52 and X63) xor (X03 and X53 and X61) xor (X03 and X53 and X63) xor (X11 and X51 and X61) xor (X11 and X51 and X62) xor (X11 and X52 and X62) xor (X11 and X52 and X63) xor (X11 and X53 and X62) xor (X12 and X51 and X62) xor (X12 and X51 and X63) xor (X12 and X52 and X61) xor (X12 and X52 and X63) xor (X12 and X53 and X61) xor (X12 and X53 and X62) xor (X13 and X51 and X62) xor (X13 and X52 and X61) xor (X13 and X52 and X63) xor (X13 and X53 and X61) xor (X13 and X53 and X63) xor (X21 and X51 and X61) xor (X21 and X51 and X62) xor (X21 and X52 and X62) xor (X21 and X52 and X63) xor (X21 and X53 and X62) xor (X22 and X51 and X62) xor (X22 and X51 and X63) xor (X22 and X52 and X61) xor (X22 and X52 and X63) xor (X22 and X53 and X61) xor (X22 and X53 and X62) xor (X23 and X51 and X62) xor (X23 and X52 and X61) xor (X23 and X52 and X63) xor (X23 and X53 and X61) xor (X23 and X53 and X63) xor (X31 and X51 and X61) xor (X31 and X51 and X62) xor (X31 and X52 and X62) xor (X31 and X52 and X63) xor (X31 and X53 and X62) xor (X32 and X51 and X62) xor (X32 and X51 and X63) xor (X32 and X52 and X61) xor (X32 and X52 and X63) xor (X32 and X53 and X61) xor (X32 and X53 and X62) xor (X33 and X51 and X62) xor (X33 and X52 and X61) xor (X33 and X52 and X63) xor (X33 and X53 and X61) xor (X33 and X53 and X63) xor (X41 and X51 and X61) xor (X41 and X51 and X62) xor (X41 and X52 and X62) xor (X41 and X52 and X63) xor (X41 and X53 and X62) xor (X42 and X51 and X62) xor (X42 and X51 and X63) xor (X42 and X52 and X61) xor (X42 and X52 and X63) xor (X42 and X53 and X61) xor (X42 and X53 and X62) xor (X43 and X51 and X62) xor (X43 and X52 and X61) xor (X43 and X52 and X63) xor (X43 and X53 and X61) xor (X43 and X53 and X63) xor (X71) xor (X0_1 and X21 and X71) xor (X0_1 and X21 and X72) xor (X0_1 and X22 and X72) xor (X0_1 and X22 and X73) xor (X0_1 and X23 and X72) xor (X02 and X21 and X72) xor (X02 and X21 and X73) xor (X02 and X22 and X71) xor (X02 and X22 and X73) xor (X02 and X23 and X71) xor (X02 and X23 and X72) xor (X03 and X21 and X72) xor (X03 and X22 and X71) xor (X03 and X22 and X73) xor (X03 and X23 and X71) xor (X03 and X23 and X73) xor (X11 and X31 and X71) xor (X11 and X31 and X72) xor (X11 and X32 and X72) xor (X11 and X32 and X73) xor (X11 and X33 and X72) xor (X12 and X31 and X72) xor (X12 and X31 and X73) xor (X12 and X32 and X71) xor (X12 and X32 and X73) xor (X12 and X33 and X71) xor (X12 and X33 and X72) xor (X13 and X31 and X72) xor (X13 and X32 and X71) xor (X13 and X32 and X73) xor (X13 and X33 and X71) xor (X13 and X33 and X73) xor (X0_1 and X41 and X71) xor (X0_1 and X41 and X72) xor (X0_1 and X42 and X72) xor (X0_1 and X42 and X73) xor (X0_1 and X43 and X72) xor (X02 and X41 and X72) xor (X02 and X41 and X73) xor (X02 and X42 and X71) xor (X02 and X42 and X73) xor (X02 and X43 and X71) xor (X02 and X43 and X72) xor (X03 and X41 and X72) xor (X03 and X42 and X71) xor (X03 and X42 and X73) xor (X03 and X43 and X71) xor (X03 and X43 and X73) xor (X51 and X71) xor (X51 and X72) xor (X52 and X71) xor (X51 and X73) xor (X0_1 and X51 and X71) xor (X0_1 and X51 and X72) xor (X0_1 and X52 and X72) xor (X0_1 and X52 and X73) xor (X0_1 and X53 and X72) xor (X02 and X51 and X72) xor (X02 and X51 and X73) xor (X02 and X52 and X71) xor (X02 and X52 and X73) xor (X02 and X53 and X71) xor (X02 and X53 and X72) xor (X03 and X51 and X72) xor (X03 and X52 and X71) xor (X03 and X52 and X73) xor (X03 and X53 and X71) xor (X03 and X53 and X73) xor (X11 and X51 and X71) xor (X11 and X51 and X72) xor (X11 and X52 and X72) xor (X11 and X52 and X73) xor (X11 and X53 and X72) xor (X12 and X51 and X72) xor (X12 and X51 and X73) xor (X12 and X52 and X71) xor (X12 and X52 and X73) xor (X12 and X53 and X71) xor (X12 and X53 and X72) xor (X13 and X51 and X72) xor (X13 and X52 and X71) xor (X13 and X52 and X73) xor (X13 and X53 and X71) xor (X13 and X53 and X73) xor (X31 and X51 and X71) xor (X31 and X51 and X72) xor (X31 and X52 and X72) xor (X31 and X52 and X73) xor (X31 and X53 and X72) xor (X32 and X51 and X72) xor (X32 and X51 and X73) xor (X32 and X52 and X71) xor (X32 and X52 and X73) xor (X32 and X53 and X71) xor (X32 and X53 and X72) xor (X33 and X51 and X72) xor (X33 and X52 and X71) xor (X33 and X52 and X73) xor (X33 and X53 and X71) xor (X33 and X53 and X73) xor (X0_1 and X61 and X71) xor (X0_1 and X61 and X72) xor (X0_1 and X62 and X72) xor (X0_1 and X62 and X73) xor (X0_1 and X63 and X72) xor (X02 and X61 and X72) xor (X02 and X61 and X73) xor (X02 and X62 and X71) xor (X02 and X62 and X73) xor (X02 and X63 and X71) xor (X02 and X63 and X72) xor (X03 and X61 and X72) xor (X03 and X62 and X71) xor (X03 and X62 and X73) xor (X03 and X63 and X71) xor (X03 and X63 and X73) xor (X21 and X61 and X71) xor (X21 and X61 and X72) xor (X21 and X62 and X72) xor (X21 and X62 and X73) xor (X21 and X63 and X72) xor (X22 and X61 and X72) xor (X22 and X61 and X73) xor (X22 and X62 and X71) xor (X22 and X62 and X73) xor (X22 and X63 and X71) xor (X22 and X63 and X72) xor (X23 and X61 and X72) xor (X23 and X62 and X71) xor (X23 and X62 and X73) xor (X23 and X63 and X71) xor (X23 and X63 and X73) xor (X41 and X61 and X71) xor (X41 and X61 and X72) xor (X41 and X62 and X72) xor (X41 and X62 and X73) xor (X41 and X63 and X72) xor (X42 and X61 and X72) xor (X42 and X61 and X73) xor (X42 and X62 and X71) xor (X42 and X62 and X73) xor (X42 and X63 and X71) xor (X42 and X63 and X72) xor (X43 and X61 and X72) xor (X43 and X62 and X71) xor (X43 and X62 and X73) xor (X43 and X63 and X71) xor (X43 and X63 and X73));
    F32  <= ((X12) xor (X02 and X12) xor (X00 and X13) xor (X02 and X13) xor (X03 and X12) xor (X12 and X22) xor (X10 and X23) xor (X12 and X23) xor (X13 and X22) xor (X00 and X10 and X23) xor (X00 and X12 and X20) xor (X00 and X12 and X22) xor (X00 and X12 and X23) xor (X00 and X13 and X20) xor (X00 and X13 and X22) xor (X02 and X10 and X22) xor (X02 and X10 and X23) xor (X02 and X13 and X20) xor (X02 and X13 and X23) xor (X03 and X10 and X20) xor (X03 and X10 and X22) xor (X03 and X10 and X23) xor (X03 and X12 and X20) xor (X03 and X12 and X22) xor (X03 and X13 and X22) xor (X32) xor (X00 and X10 and X33) xor (X00 and X12 and X30) xor (X00 and X12 and X32) xor (X00 and X12 and X33) xor (X00 and X13 and X30) xor (X00 and X13 and X32) xor (X02 and X10 and X32) xor (X02 and X10 and X33) xor (X02 and X13 and X30) xor (X02 and X13 and X33) xor (X03 and X10 and X30) xor (X03 and X10 and X32) xor (X03 and X10 and X33) xor (X03 and X12 and X30) xor (X03 and X12 and X32) xor (X03 and X13 and X32) xor (X22 and X32) xor (X20 and X33) xor (X22 and X33) xor (X23 and X32) xor (X42) xor (X02 and X42) xor (X00 and X43) xor (X02 and X43) xor (X03 and X42) xor (X00 and X10 and X43) xor (X00 and X12 and X40) xor (X00 and X12 and X42) xor (X00 and X12 and X43) xor (X00 and X13 and X40) xor (X00 and X13 and X42) xor (X02 and X10 and X42) xor (X02 and X10 and X43) xor (X02 and X13 and X40) xor (X02 and X13 and X43) xor (X03 and X10 and X40) xor (X03 and X10 and X42) xor (X03 and X10 and X43) xor (X03 and X12 and X40) xor (X03 and X12 and X42) xor (X03 and X13 and X42) xor (X22 and X42) xor (X20 and X43) xor (X22 and X43) xor (X23 and X42) xor (X00 and X20 and X43) xor (X00 and X22 and X40) xor (X00 and X22 and X42) xor (X00 and X22 and X43) xor (X00 and X23 and X40) xor (X00 and X23 and X42) xor (X02 and X20 and X42) xor (X02 and X20 and X43) xor (X02 and X23 and X40) xor (X02 and X23 and X43) xor (X03 and X20 and X40) xor (X03 and X20 and X42) xor (X03 and X20 and X43) xor (X03 and X22 and X40) xor (X03 and X22 and X42) xor (X03 and X23 and X42) xor (X10 and X20 and X43) xor (X10 and X22 and X40) xor (X10 and X22 and X42) xor (X10 and X22 and X43) xor (X10 and X23 and X40) xor (X10 and X23 and X42) xor (X12 and X20 and X42) xor (X12 and X20 and X43) xor (X12 and X23 and X40) xor (X12 and X23 and X43) xor (X13 and X20 and X40) xor (X13 and X20 and X42) xor (X13 and X20 and X43) xor (X13 and X22 and X40) xor (X13 and X22 and X42) xor (X13 and X23 and X42) xor (X32 and X42) xor (X30 and X43) xor (X32 and X43) xor (X33 and X42) xor (X12 and X52) xor (X10 and X53) xor (X12 and X53) xor (X13 and X52) xor (X22 and X52) xor (X20 and X53) xor (X22 and X53) xor (X23 and X52) xor (X20 and X30 and X53) xor (X20 and X32 and X50) xor (X20 and X32 and X52) xor (X20 and X32 and X53) xor (X20 and X33 and X50) xor (X20 and X33 and X52) xor (X22 and X30 and X52) xor (X22 and X30 and X53) xor (X22 and X33 and X50) xor (X22 and X33 and X53) xor (X23 and X30 and X50) xor (X23 and X30 and X52) xor (X23 and X30 and X53) xor (X23 and X32 and X50) xor (X23 and X32 and X52) xor (X23 and X33 and X52) xor (X00 and X40 and X53) xor (X00 and X42 and X50) xor (X00 and X42 and X52) xor (X00 and X42 and X53) xor (X00 and X43 and X50) xor (X00 and X43 and X52) xor (X02 and X40 and X52) xor (X02 and X40 and X53) xor (X02 and X43 and X50) xor (X02 and X43 and X53) xor (X03 and X40 and X50) xor (X03 and X40 and X52) xor (X03 and X40 and X53) xor (X03 and X42 and X50) xor (X03 and X42 and X52) xor (X03 and X43 and X52) xor (X10 and X40 and X53) xor (X10 and X42 and X50) xor (X10 and X42 and X52) xor (X10 and X42 and X53) xor (X10 and X43 and X50) xor (X10 and X43 and X52) xor (X12 and X40 and X52) xor (X12 and X40 and X53) xor (X12 and X43 and X50) xor (X12 and X43 and X53) xor (X13 and X40 and X50) xor (X13 and X40 and X52) xor (X13 and X40 and X53) xor (X13 and X42 and X50) xor (X13 and X42 and X52) xor (X13 and X43 and X52) xor (X30 and X40 and X53) xor (X30 and X42 and X50) xor (X30 and X42 and X52) xor (X30 and X42 and X53) xor (X30 and X43 and X50) xor (X30 and X43 and X52) xor (X32 and X40 and X52) xor (X32 and X40 and X53) xor (X32 and X43 and X50) xor (X32 and X43 and X53) xor (X33 and X40 and X50) xor (X33 and X40 and X52) xor (X33 and X40 and X53) xor (X33 and X42 and X50) xor (X33 and X42 and X52) xor (X33 and X43 and X52) xor (X62) xor (X02 and X62) xor (X00 and X63) xor (X02 and X63) xor (X03 and X62) xor (X00 and X10 and X63) xor (X00 and X12 and X60) xor (X00 and X12 and X62) xor (X00 and X12 and X63) xor (X00 and X13 and X60) xor (X00 and X13 and X62) xor (X02 and X10 and X62) xor (X02 and X10 and X63) xor (X02 and X13 and X60) xor (X02 and X13 and X63) xor (X03 and X10 and X60) xor (X03 and X10 and X62) xor (X03 and X10 and X63) xor (X03 and X12 and X60) xor (X03 and X12 and X62) xor (X03 and X13 and X62) xor (X22 and X62) xor (X20 and X63) xor (X22 and X63) xor (X23 and X62) xor (X10 and X20 and X63) xor (X10 and X22 and X60) xor (X10 and X22 and X62) xor (X10 and X22 and X63) xor (X10 and X23 and X60) xor (X10 and X23 and X62) xor (X12 and X20 and X62) xor (X12 and X20 and X63) xor (X12 and X23 and X60) xor (X12 and X23 and X63) xor (X13 and X20 and X60) xor (X13 and X20 and X62) xor (X13 and X20 and X63) xor (X13 and X22 and X60) xor (X13 and X22 and X62) xor (X13 and X23 and X62) xor (X32 and X62) xor (X30 and X63) xor (X32 and X63) xor (X33 and X62) xor (X00 and X30 and X63) xor (X00 and X32 and X60) xor (X00 and X32 and X62) xor (X00 and X32 and X63) xor (X00 and X33 and X60) xor (X00 and X33 and X62) xor (X02 and X30 and X62) xor (X02 and X30 and X63) xor (X02 and X33 and X60) xor (X02 and X33 and X63) xor (X03 and X30 and X60) xor (X03 and X30 and X62) xor (X03 and X30 and X63) xor (X03 and X32 and X60) xor (X03 and X32 and X62) xor (X03 and X33 and X62) xor (X42 and X62) xor (X40 and X63) xor (X42 and X63) xor (X43 and X62) xor (X10 and X40 and X63) xor (X10 and X42 and X60) xor (X10 and X42 and X62) xor (X10 and X42 and X63) xor (X10 and X43 and X60) xor (X10 and X43 and X62) xor (X12 and X40 and X62) xor (X12 and X40 and X63) xor (X12 and X43 and X60) xor (X12 and X43 and X63) xor (X13 and X40 and X60) xor (X13 and X40 and X62) xor (X13 and X40 and X63) xor (X13 and X42 and X60) xor (X13 and X42 and X62) xor (X13 and X43 and X62) xor (X52 and X62) xor (X50 and X63) xor (X52 and X63) xor (X53 and X62) xor (X00 and X50 and X63) xor (X00 and X52 and X60) xor (X00 and X52 and X62) xor (X00 and X52 and X63) xor (X00 and X53 and X60) xor (X00 and X53 and X62) xor (X02 and X50 and X62) xor (X02 and X50 and X63) xor (X02 and X53 and X60) xor (X02 and X53 and X63) xor (X03 and X50 and X60) xor (X03 and X50 and X62) xor (X03 and X50 and X63) xor (X03 and X52 and X60) xor (X03 and X52 and X62) xor (X03 and X53 and X62) xor (X10 and X50 and X63) xor (X10 and X52 and X60) xor (X10 and X52 and X62) xor (X10 and X52 and X63) xor (X10 and X53 and X60) xor (X10 and X53 and X62) xor (X12 and X50 and X62) xor (X12 and X50 and X63) xor (X12 and X53 and X60) xor (X12 and X53 and X63) xor (X13 and X50 and X60) xor (X13 and X50 and X62) xor (X13 and X50 and X63) xor (X13 and X52 and X60) xor (X13 and X52 and X62) xor (X13 and X53 and X62) xor (X20 and X50 and X63) xor (X20 and X52 and X60) xor (X20 and X52 and X62) xor (X20 and X52 and X63) xor (X20 and X53 and X60) xor (X20 and X53 and X62) xor (X22 and X50 and X62) xor (X22 and X50 and X63) xor (X22 and X53 and X60) xor (X22 and X53 and X63) xor (X23 and X50 and X60) xor (X23 and X50 and X62) xor (X23 and X50 and X63) xor (X23 and X52 and X60) xor (X23 and X52 and X62) xor (X23 and X53 and X62) xor (X30 and X50 and X63) xor (X30 and X52 and X60) xor (X30 and X52 and X62) xor (X30 and X52 and X63) xor (X30 and X53 and X60) xor (X30 and X53 and X62) xor (X32 and X50 and X62) xor (X32 and X50 and X63) xor (X32 and X53 and X60) xor (X32 and X53 and X63) xor (X33 and X50 and X60) xor (X33 and X50 and X62) xor (X33 and X50 and X63) xor (X33 and X52 and X60) xor (X33 and X52 and X62) xor (X33 and X53 and X62) xor (X40 and X50 and X63) xor (X40 and X52 and X60) xor (X40 and X52 and X62) xor (X40 and X52 and X63) xor (X40 and X53 and X60) xor (X40 and X53 and X62) xor (X42 and X50 and X62) xor (X42 and X50 and X63) xor (X42 and X53 and X60) xor (X42 and X53 and X63) xor (X43 and X50 and X60) xor (X43 and X50 and X62) xor (X43 and X50 and X63) xor (X43 and X52 and X60) xor (X43 and X52 and X62) xor (X43 and X53 and X62) xor (X72) xor (X00 and X20 and X73) xor (X00 and X22 and X70) xor (X00 and X22 and X72) xor (X00 and X22 and X73) xor (X00 and X23 and X70) xor (X00 and X23 and X72) xor (X02 and X20 and X72) xor (X02 and X20 and X73) xor (X02 and X23 and X70) xor (X02 and X23 and X73) xor (X03 and X20 and X70) xor (X03 and X20 and X72) xor (X03 and X20 and X73) xor (X03 and X22 and X70) xor (X03 and X22 and X72) xor (X03 and X23 and X72) xor (X10 and X30 and X73) xor (X10 and X32 and X70) xor (X10 and X32 and X72) xor (X10 and X32 and X73) xor (X10 and X33 and X70) xor (X10 and X33 and X72) xor (X12 and X30 and X72) xor (X12 and X30 and X73) xor (X12 and X33 and X70) xor (X12 and X33 and X73) xor (X13 and X30 and X70) xor (X13 and X30 and X72) xor (X13 and X30 and X73) xor (X13 and X32 and X70) xor (X13 and X32 and X72) xor (X13 and X33 and X72) xor (X00 and X40 and X73) xor (X00 and X42 and X70) xor (X00 and X42 and X72) xor (X00 and X42 and X73) xor (X00 and X43 and X70) xor (X00 and X43 and X72) xor (X02 and X40 and X72) xor (X02 and X40 and X73) xor (X02 and X43 and X70) xor (X02 and X43 and X73) xor (X03 and X40 and X70) xor (X03 and X40 and X72) xor (X03 and X40 and X73) xor (X03 and X42 and X70) xor (X03 and X42 and X72) xor (X03 and X43 and X72) xor (X52 and X72) xor (X50 and X73) xor (X52 and X73) xor (X53 and X72) xor (X00 and X50 and X73) xor (X00 and X52 and X70) xor (X00 and X52 and X72) xor (X00 and X52 and X73) xor (X00 and X53 and X70) xor (X00 and X53 and X72) xor (X02 and X50 and X72) xor (X02 and X50 and X73) xor (X02 and X53 and X70) xor (X02 and X53 and X73) xor (X03 and X50 and X70) xor (X03 and X50 and X72) xor (X03 and X50 and X73) xor (X03 and X52 and X70) xor (X03 and X52 and X72) xor (X03 and X53 and X72) xor (X10 and X50 and X73) xor (X10 and X52 and X70) xor (X10 and X52 and X72) xor (X10 and X52 and X73) xor (X10 and X53 and X70) xor (X10 and X53 and X72) xor (X12 and X50 and X72) xor (X12 and X50 and X73) xor (X12 and X53 and X70) xor (X12 and X53 and X73) xor (X13 and X50 and X70) xor (X13 and X50 and X72) xor (X13 and X50 and X73) xor (X13 and X52 and X70) xor (X13 and X52 and X72) xor (X13 and X53 and X72) xor (X30 and X50 and X73) xor (X30 and X52 and X70) xor (X30 and X52 and X72) xor (X30 and X52 and X73) xor (X30 and X53 and X70) xor (X30 and X53 and X72) xor (X32 and X50 and X72) xor (X32 and X50 and X73) xor (X32 and X53 and X70) xor (X32 and X53 and X73) xor (X33 and X50 and X70) xor (X33 and X50 and X72) xor (X33 and X50 and X73) xor (X33 and X52 and X70) xor (X33 and X52 and X72) xor (X33 and X53 and X72) xor (X00 and X60 and X73) xor (X00 and X62 and X70) xor (X00 and X62 and X72) xor (X00 and X62 and X73) xor (X00 and X63 and X70) xor (X00 and X63 and X72) xor (X02 and X60 and X72) xor (X02 and X60 and X73) xor (X02 and X63 and X70) xor (X02 and X63 and X73) xor (X03 and X60 and X70) xor (X03 and X60 and X72) xor (X03 and X60 and X73) xor (X03 and X62 and X70) xor (X03 and X62 and X72) xor (X03 and X63 and X72) xor (X20 and X60 and X73) xor (X20 and X62 and X70) xor (X20 and X62 and X72) xor (X20 and X62 and X73) xor (X20 and X63 and X70) xor (X20 and X63 and X72) xor (X22 and X60 and X72) xor (X22 and X60 and X73) xor (X22 and X63 and X70) xor (X22 and X63 and X73) xor (X23 and X60 and X70) xor (X23 and X60 and X72) xor (X23 and X60 and X73) xor (X23 and X62 and X70) xor (X23 and X62 and X72) xor (X23 and X63 and X72) xor (X40 and X60 and X73) xor (X40 and X62 and X70) xor (X40 and X62 and X72) xor (X40 and X62 and X73) xor (X40 and X63 and X70) xor (X40 and X63 and X72) xor (X42 and X60 and X72) xor (X42 and X60 and X73) xor (X42 and X63 and X70) xor (X42 and X63 and X73) xor (X43 and X60 and X70) xor (X43 and X60 and X72) xor (X43 and X60 and X73) xor (X43 and X62 and X70) xor (X43 and X62 and X72) xor (X43 and X63 and X72));
    F33  <= ((X13) xor (X03 and X13) xor (X03 and X10) xor (X03 and X11) xor (X0_1 and X10) xor (X13 and X23) xor (X13 and X20) xor (X13 and X21) xor (X11 and X20) xor (X00 and X10 and X21) xor (X00 and X11 and X20) xor (X00 and X11 and X23) xor (X00 and X13 and X21) xor (X00 and X13 and X23) xor (X0_1 and X10 and X21) xor (X0_1 and X10 and X23) xor (X0_1 and X11 and X23) xor (X0_1 and X13 and X20) xor (X0_1 and X13 and X21) xor (X0_1 and X13 and X23) xor (X03 and X10 and X21) xor (X03 and X11 and X20) xor (X03 and X11 and X21) xor (X03 and X11 and X23) xor (X03 and X13 and X20) xor (X33) xor (X00 and X10 and X31) xor (X00 and X11 and X30) xor (X00 and X11 and X33) xor (X00 and X13 and X31) xor (X00 and X13 and X33) xor (X0_1 and X10 and X31) xor (X0_1 and X10 and X33) xor (X0_1 and X11 and X33) xor (X0_1 and X13 and X30) xor (X0_1 and X13 and X31) xor (X0_1 and X13 and X33) xor (X03 and X10 and X31) xor (X03 and X11 and X30) xor (X03 and X11 and X31) xor (X03 and X11 and X33) xor (X03 and X13 and X30) xor (X23 and X33) xor (X23 and X30) xor (X23 and X31) xor (X21 and X30) xor (X43) xor (X03 and X43) xor (X03 and X40) xor (X03 and X41) xor (X0_1 and X40) xor (X00 and X10 and X41) xor (X00 and X11 and X40) xor (X00 and X11 and X43) xor (X00 and X13 and X41) xor (X00 and X13 and X43) xor (X0_1 and X10 and X41) xor (X0_1 and X10 and X43) xor (X0_1 and X11 and X43) xor (X0_1 and X13 and X40) xor (X0_1 and X13 and X41) xor (X0_1 and X13 and X43) xor (X03 and X10 and X41) xor (X03 and X11 and X40) xor (X03 and X11 and X41) xor (X03 and X11 and X43) xor (X03 and X13 and X40) xor (X23 and X43) xor (X23 and X40) xor (X23 and X41) xor (X21 and X40) xor (X00 and X20 and X41) xor (X00 and X21 and X40) xor (X00 and X21 and X43) xor (X00 and X23 and X41) xor (X00 and X23 and X43) xor (X0_1 and X20 and X41) xor (X0_1 and X20 and X43) xor (X0_1 and X21 and X43) xor (X0_1 and X23 and X40) xor (X0_1 and X23 and X41) xor (X0_1 and X23 and X43) xor (X03 and X20 and X41) xor (X03 and X21 and X40) xor (X03 and X21 and X41) xor (X03 and X21 and X43) xor (X03 and X23 and X40) xor (X10 and X20 and X41) xor (X10 and X21 and X40) xor (X10 and X21 and X43) xor (X10 and X23 and X41) xor (X10 and X23 and X43) xor (X11 and X20 and X41) xor (X11 and X20 and X43) xor (X11 and X21 and X43) xor (X11 and X23 and X40) xor (X11 and X23 and X41) xor (X11 and X23 and X43) xor (X13 and X20 and X41) xor (X13 and X21 and X40) xor (X13 and X21 and X41) xor (X13 and X21 and X43) xor (X13 and X23 and X40) xor (X33 and X43) xor (X33 and X40) xor (X33 and X41) xor (X31 and X40) xor (X13 and X53) xor (X13 and X50) xor (X13 and X51) xor (X11 and X50) xor (X23 and X53) xor (X23 and X50) xor (X23 and X51) xor (X21 and X50) xor (X20 and X30 and X51) xor (X20 and X31 and X50) xor (X20 and X31 and X53) xor (X20 and X33 and X51) xor (X20 and X33 and X53) xor (X21 and X30 and X51) xor (X21 and X30 and X53) xor (X21 and X31 and X53) xor (X21 and X33 and X50) xor (X21 and X33 and X51) xor (X21 and X33 and X53) xor (X23 and X30 and X51) xor (X23 and X31 and X50) xor (X23 and X31 and X51) xor (X23 and X31 and X53) xor (X23 and X33 and X50) xor (X00 and X40 and X51) xor (X00 and X41 and X50) xor (X00 and X41 and X53) xor (X00 and X43 and X51) xor (X00 and X43 and X53) xor (X0_1 and X40 and X51) xor (X0_1 and X40 and X53) xor (X0_1 and X41 and X53) xor (X0_1 and X43 and X50) xor (X0_1 and X43 and X51) xor (X0_1 and X43 and X53) xor (X03 and X40 and X51) xor (X03 and X41 and X50) xor (X03 and X41 and X51) xor (X03 and X41 and X53) xor (X03 and X43 and X50) xor (X10 and X40 and X51) xor (X10 and X41 and X50) xor (X10 and X41 and X53) xor (X10 and X43 and X51) xor (X10 and X43 and X53) xor (X11 and X40 and X51) xor (X11 and X40 and X53) xor (X11 and X41 and X53) xor (X11 and X43 and X50) xor (X11 and X43 and X51) xor (X11 and X43 and X53) xor (X13 and X40 and X51) xor (X13 and X41 and X50) xor (X13 and X41 and X51) xor (X13 and X41 and X53) xor (X13 and X43 and X50) xor (X30 and X40 and X51) xor (X30 and X41 and X50) xor (X30 and X41 and X53) xor (X30 and X43 and X51) xor (X30 and X43 and X53) xor (X31 and X40 and X51) xor (X31 and X40 and X53) xor (X31 and X41 and X53) xor (X31 and X43 and X50) xor (X31 and X43 and X51) xor (X31 and X43 and X53) xor (X33 and X40 and X51) xor (X33 and X41 and X50) xor (X33 and X41 and X51) xor (X33 and X41 and X53) xor (X33 and X43 and X50) xor (X63) xor (X03 and X63) xor (X03 and X60) xor (X03 and X61) xor (X0_1 and X60) xor (X00 and X10 and X61) xor (X00 and X11 and X60) xor (X00 and X11 and X63) xor (X00 and X13 and X61) xor (X00 and X13 and X63) xor (X0_1 and X10 and X61) xor (X0_1 and X10 and X63) xor (X0_1 and X11 and X63) xor (X0_1 and X13 and X60) xor (X0_1 and X13 and X61) xor (X0_1 and X13 and X63) xor (X03 and X10 and X61) xor (X03 and X11 and X60) xor (X03 and X11 and X61) xor (X03 and X11 and X63) xor (X03 and X13 and X60) xor (X23 and X63) xor (X23 and X60) xor (X23 and X61) xor (X21 and X60) xor (X10 and X20 and X61) xor (X10 and X21 and X60) xor (X10 and X21 and X63) xor (X10 and X23 and X61) xor (X10 and X23 and X63) xor (X11 and X20 and X61) xor (X11 and X20 and X63) xor (X11 and X21 and X63) xor (X11 and X23 and X60) xor (X11 and X23 and X61) xor (X11 and X23 and X63) xor (X13 and X20 and X61) xor (X13 and X21 and X60) xor (X13 and X21 and X61) xor (X13 and X21 and X63) xor (X13 and X23 and X60) xor (X33 and X63) xor (X33 and X60) xor (X33 and X61) xor (X31 and X60) xor (X00 and X30 and X61) xor (X00 and X31 and X60) xor (X00 and X31 and X63) xor (X00 and X33 and X61) xor (X00 and X33 and X63) xor (X0_1 and X30 and X61) xor (X0_1 and X30 and X63) xor (X0_1 and X31 and X63) xor (X0_1 and X33 and X60) xor (X0_1 and X33 and X61) xor (X0_1 and X33 and X63) xor (X03 and X30 and X61) xor (X03 and X31 and X60) xor (X03 and X31 and X61) xor (X03 and X31 and X63) xor (X03 and X33 and X60) xor (X43 and X63) xor (X43 and X60) xor (X43 and X61) xor (X41 and X60) xor (X10 and X40 and X61) xor (X10 and X41 and X60) xor (X10 and X41 and X63) xor (X10 and X43 and X61) xor (X10 and X43 and X63) xor (X11 and X40 and X61) xor (X11 and X40 and X63) xor (X11 and X41 and X63) xor (X11 and X43 and X60) xor (X11 and X43 and X61) xor (X11 and X43 and X63) xor (X13 and X40 and X61) xor (X13 and X41 and X60) xor (X13 and X41 and X61) xor (X13 and X41 and X63) xor (X13 and X43 and X60) xor (X53 and X63) xor (X53 and X60) xor (X53 and X61) xor (X51 and X60) xor (X00 and X50 and X61) xor (X00 and X51 and X60) xor (X00 and X51 and X63) xor (X00 and X53 and X61) xor (X00 and X53 and X63) xor (X0_1 and X50 and X61) xor (X0_1 and X50 and X63) xor (X0_1 and X51 and X63) xor (X0_1 and X53 and X60) xor (X0_1 and X53 and X61) xor (X0_1 and X53 and X63) xor (X03 and X50 and X61) xor (X03 and X51 and X60) xor (X03 and X51 and X61) xor (X03 and X51 and X63) xor (X03 and X53 and X60) xor (X10 and X50 and X61) xor (X10 and X51 and X60) xor (X10 and X51 and X63) xor (X10 and X53 and X61) xor (X10 and X53 and X63) xor (X11 and X50 and X61) xor (X11 and X50 and X63) xor (X11 and X51 and X63) xor (X11 and X53 and X60) xor (X11 and X53 and X61) xor (X11 and X53 and X63) xor (X13 and X50 and X61) xor (X13 and X51 and X60) xor (X13 and X51 and X61) xor (X13 and X51 and X63) xor (X13 and X53 and X60) xor (X20 and X50 and X61) xor (X20 and X51 and X60) xor (X20 and X51 and X63) xor (X20 and X53 and X61) xor (X20 and X53 and X63) xor (X21 and X50 and X61) xor (X21 and X50 and X63) xor (X21 and X51 and X63) xor (X21 and X53 and X60) xor (X21 and X53 and X61) xor (X21 and X53 and X63) xor (X23 and X50 and X61) xor (X23 and X51 and X60) xor (X23 and X51 and X61) xor (X23 and X51 and X63) xor (X23 and X53 and X60) xor (X30 and X50 and X61) xor (X30 and X51 and X60) xor (X30 and X51 and X63) xor (X30 and X53 and X61) xor (X30 and X53 and X63) xor (X31 and X50 and X61) xor (X31 and X50 and X63) xor (X31 and X51 and X63) xor (X31 and X53 and X60) xor (X31 and X53 and X61) xor (X31 and X53 and X63) xor (X33 and X50 and X61) xor (X33 and X51 and X60) xor (X33 and X51 and X61) xor (X33 and X51 and X63) xor (X33 and X53 and X60) xor (X40 and X50 and X61) xor (X40 and X51 and X60) xor (X40 and X51 and X63) xor (X40 and X53 and X61) xor (X40 and X53 and X63) xor (X41 and X50 and X61) xor (X41 and X50 and X63) xor (X41 and X51 and X63) xor (X41 and X53 and X60) xor (X41 and X53 and X61) xor (X41 and X53 and X63) xor (X43 and X50 and X61) xor (X43 and X51 and X60) xor (X43 and X51 and X61) xor (X43 and X51 and X63) xor (X43 and X53 and X60) xor (X73) xor (X00 and X20 and X71) xor (X00 and X21 and X70) xor (X00 and X21 and X73) xor (X00 and X23 and X71) xor (X00 and X23 and X73) xor (X0_1 and X20 and X71) xor (X0_1 and X20 and X73) xor (X0_1 and X21 and X73) xor (X0_1 and X23 and X70) xor (X0_1 and X23 and X71) xor (X0_1 and X23 and X73) xor (X03 and X20 and X71) xor (X03 and X21 and X70) xor (X03 and X21 and X71) xor (X03 and X21 and X73) xor (X03 and X23 and X70) xor (X10 and X30 and X71) xor (X10 and X31 and X70) xor (X10 and X31 and X73) xor (X10 and X33 and X71) xor (X10 and X33 and X73) xor (X11 and X30 and X71) xor (X11 and X30 and X73) xor (X11 and X31 and X73) xor (X11 and X33 and X70) xor (X11 and X33 and X71) xor (X11 and X33 and X73) xor (X13 and X30 and X71) xor (X13 and X31 and X70) xor (X13 and X31 and X71) xor (X13 and X31 and X73) xor (X13 and X33 and X70) xor (X00 and X40 and X71) xor (X00 and X41 and X70) xor (X00 and X41 and X73) xor (X00 and X43 and X71) xor (X00 and X43 and X73) xor (X0_1 and X40 and X71) xor (X0_1 and X40 and X73) xor (X0_1 and X41 and X73) xor (X0_1 and X43 and X70) xor (X0_1 and X43 and X71) xor (X0_1 and X43 and X73) xor (X03 and X40 and X71) xor (X03 and X41 and X70) xor (X03 and X41 and X71) xor (X03 and X41 and X73) xor (X03 and X43 and X70) xor (X53 and X73) xor (X53 and X70) xor (X53 and X71) xor (X51 and X70) xor (X00 and X50 and X71) xor (X00 and X51 and X70) xor (X00 and X51 and X73) xor (X00 and X53 and X71) xor (X00 and X53 and X73) xor (X0_1 and X50 and X71) xor (X0_1 and X50 and X73) xor (X0_1 and X51 and X73) xor (X0_1 and X53 and X70) xor (X0_1 and X53 and X71) xor (X0_1 and X53 and X73) xor (X03 and X50 and X71) xor (X03 and X51 and X70) xor (X03 and X51 and X71) xor (X03 and X51 and X73) xor (X03 and X53 and X70) xor (X10 and X50 and X71) xor (X10 and X51 and X70) xor (X10 and X51 and X73) xor (X10 and X53 and X71) xor (X10 and X53 and X73) xor (X11 and X50 and X71) xor (X11 and X50 and X73) xor (X11 and X51 and X73) xor (X11 and X53 and X70) xor (X11 and X53 and X71) xor (X11 and X53 and X73) xor (X13 and X50 and X71) xor (X13 and X51 and X70) xor (X13 and X51 and X71) xor (X13 and X51 and X73) xor (X13 and X53 and X70) xor (X30 and X50 and X71) xor (X30 and X51 and X70) xor (X30 and X51 and X73) xor (X30 and X53 and X71) xor (X30 and X53 and X73) xor (X31 and X50 and X71) xor (X31 and X50 and X73) xor (X31 and X51 and X73) xor (X31 and X53 and X70) xor (X31 and X53 and X71) xor (X31 and X53 and X73) xor (X33 and X50 and X71) xor (X33 and X51 and X70) xor (X33 and X51 and X71) xor (X33 and X51 and X73) xor (X33 and X53 and X70) xor (X00 and X60 and X71) xor (X00 and X61 and X70) xor (X00 and X61 and X73) xor (X00 and X63 and X71) xor (X00 and X63 and X73) xor (X0_1 and X60 and X71) xor (X0_1 and X60 and X73) xor (X0_1 and X61 and X73) xor (X0_1 and X63 and X70) xor (X0_1 and X63 and X71) xor (X0_1 and X63 and X73) xor (X03 and X60 and X71) xor (X03 and X61 and X70) xor (X03 and X61 and X71) xor (X03 and X61 and X73) xor (X03 and X63 and X70) xor (X20 and X60 and X71) xor (X20 and X61 and X70) xor (X20 and X61 and X73) xor (X20 and X63 and X71) xor (X20 and X63 and X73) xor (X21 and X60 and X71) xor (X21 and X60 and X73) xor (X21 and X61 and X73) xor (X21 and X63 and X70) xor (X21 and X63 and X71) xor (X21 and X63 and X73) xor (X23 and X60 and X71) xor (X23 and X61 and X70) xor (X23 and X61 and X71) xor (X23 and X61 and X73) xor (X23 and X63 and X70) xor (X40 and X60 and X71) xor (X40 and X61 and X70) xor (X40 and X61 and X73) xor (X40 and X63 and X71) xor (X40 and X63 and X73) xor (X41 and X60 and X71) xor (X41 and X60 and X73) xor (X41 and X61 and X73) xor (X41 and X63 and X70) xor (X41 and X63 and X71) xor (X41 and X63 and X73) xor (X43 and X60 and X71) xor (X43 and X61 and X70) xor (X43 and X61 and X71) xor (X43 and X61 and X73) xor (X43 and X63 and X70));
    F40  <= ((X00 and X10) xor (X00 and X11) xor (X02 and X10) xor (X00 and X12) xor (X20) xor (X30) xor (X00 and X30) xor (X00 and X31) xor (X02 and X30) xor (X00 and X32) xor (X20 and X30) xor (X20 and X31) xor (X22 and X30) xor (X20 and X32) xor (X00 and X20 and X30) xor (X00 and X20 and X32) xor (X00 and X21 and X31) xor (X00 and X21 and X32) xor (X00 and X22 and X31) xor (X0_1 and X20 and X30) xor (X0_1 and X20 and X32) xor (X0_1 and X21 and X30) xor (X0_1 and X22 and X30) xor (X0_1 and X22 and X31) xor (X02 and X20 and X30) xor (X02 and X20 and X31) xor (X02 and X21 and X30) xor (X02 and X21 and X31) xor (X02 and X22 and X30) xor (X02 and X22 and X32) xor (X10 and X20 and X30) xor (X10 and X20 and X32) xor (X10 and X21 and X31) xor (X10 and X21 and X32) xor (X10 and X22 and X31) xor (X11 and X20 and X30) xor (X11 and X20 and X32) xor (X11 and X21 and X30) xor (X11 and X22 and X30) xor (X11 and X22 and X31) xor (X12 and X20 and X30) xor (X12 and X20 and X31) xor (X12 and X21 and X30) xor (X12 and X21 and X31) xor (X12 and X22 and X30) xor (X12 and X22 and X32) xor (X10 and X40) xor (X10 and X41) xor (X12 and X40) xor (X10 and X42) xor (X00 and X10 and X40) xor (X00 and X10 and X42) xor (X00 and X11 and X41) xor (X00 and X11 and X42) xor (X00 and X12 and X41) xor (X0_1 and X10 and X40) xor (X0_1 and X10 and X42) xor (X0_1 and X11 and X40) xor (X0_1 and X12 and X40) xor (X0_1 and X12 and X41) xor (X02 and X10 and X40) xor (X02 and X10 and X41) xor (X02 and X11 and X40) xor (X02 and X11 and X41) xor (X02 and X12 and X40) xor (X02 and X12 and X42) xor (X30 and X40) xor (X30 and X41) xor (X32 and X40) xor (X30 and X42) xor (X00 and X30 and X40) xor (X00 and X30 and X42) xor (X00 and X31 and X41) xor (X00 and X31 and X42) xor (X00 and X32 and X41) xor (X0_1 and X30 and X40) xor (X0_1 and X30 and X42) xor (X0_1 and X31 and X40) xor (X0_1 and X32 and X40) xor (X0_1 and X32 and X41) xor (X02 and X30 and X40) xor (X02 and X30 and X41) xor (X02 and X31 and X40) xor (X02 and X31 and X41) xor (X02 and X32 and X40) xor (X02 and X32 and X42) xor (X10 and X30 and X40) xor (X10 and X30 and X42) xor (X10 and X31 and X41) xor (X10 and X31 and X42) xor (X10 and X32 and X41) xor (X11 and X30 and X40) xor (X11 and X30 and X42) xor (X11 and X31 and X40) xor (X11 and X32 and X40) xor (X11 and X32 and X41) xor (X12 and X30 and X40) xor (X12 and X30 and X41) xor (X12 and X31 and X40) xor (X12 and X31 and X41) xor (X12 and X32 and X40) xor (X12 and X32 and X42) xor (X20 and X30 and X40) xor (X20 and X30 and X42) xor (X20 and X31 and X41) xor (X20 and X31 and X42) xor (X20 and X32 and X41) xor (X21 and X30 and X40) xor (X21 and X30 and X42) xor (X21 and X31 and X40) xor (X21 and X32 and X40) xor (X21 and X32 and X41) xor (X22 and X30 and X40) xor (X22 and X30 and X41) xor (X22 and X31 and X40) xor (X22 and X31 and X41) xor (X22 and X32 and X40) xor (X22 and X32 and X42) xor (X50) xor (X10 and X50) xor (X10 and X51) xor (X12 and X50) xor (X10 and X52) xor (X00 and X10 and X50) xor (X00 and X10 and X52) xor (X00 and X11 and X51) xor (X00 and X11 and X52) xor (X00 and X12 and X51) xor (X0_1 and X10 and X50) xor (X0_1 and X10 and X52) xor (X0_1 and X11 and X50) xor (X0_1 and X12 and X50) xor (X0_1 and X12 and X51) xor (X02 and X10 and X50) xor (X02 and X10 and X51) xor (X02 and X11 and X50) xor (X02 and X11 and X51) xor (X02 and X12 and X50) xor (X02 and X12 and X52) xor (X00 and X20 and X50) xor (X00 and X20 and X52) xor (X00 and X21 and X51) xor (X00 and X21 and X52) xor (X00 and X22 and X51) xor (X0_1 and X20 and X50) xor (X0_1 and X20 and X52) xor (X0_1 and X21 and X50) xor (X0_1 and X22 and X50) xor (X0_1 and X22 and X51) xor (X02 and X20 and X50) xor (X02 and X20 and X51) xor (X02 and X21 and X50) xor (X02 and X21 and X51) xor (X02 and X22 and X50) xor (X02 and X22 and X52) xor (X10 and X20 and X50) xor (X10 and X20 and X52) xor (X10 and X21 and X51) xor (X10 and X21 and X52) xor (X10 and X22 and X51) xor (X11 and X20 and X50) xor (X11 and X20 and X52) xor (X11 and X21 and X50) xor (X11 and X22 and X50) xor (X11 and X22 and X51) xor (X12 and X20 and X50) xor (X12 and X20 and X51) xor (X12 and X21 and X50) xor (X12 and X21 and X51) xor (X12 and X22 and X50) xor (X12 and X22 and X52) xor (X30 and X50) xor (X30 and X51) xor (X32 and X50) xor (X30 and X52) xor (X10 and X30 and X50) xor (X10 and X30 and X52) xor (X10 and X31 and X51) xor (X10 and X31 and X52) xor (X10 and X32 and X51) xor (X11 and X30 and X50) xor (X11 and X30 and X52) xor (X11 and X31 and X50) xor (X11 and X32 and X50) xor (X11 and X32 and X51) xor (X12 and X30 and X50) xor (X12 and X30 and X51) xor (X12 and X31 and X50) xor (X12 and X31 and X51) xor (X12 and X32 and X50) xor (X12 and X32 and X52) xor (X20 and X30 and X50) xor (X20 and X30 and X52) xor (X20 and X31 and X51) xor (X20 and X31 and X52) xor (X20 and X32 and X51) xor (X21 and X30 and X50) xor (X21 and X30 and X52) xor (X21 and X31 and X50) xor (X21 and X32 and X50) xor (X21 and X32 and X51) xor (X22 and X30 and X50) xor (X22 and X30 and X51) xor (X22 and X31 and X50) xor (X22 and X31 and X51) xor (X22 and X32 and X50) xor (X22 and X32 and X52) xor (X40 and X50) xor (X40 and X51) xor (X42 and X50) xor (X40 and X52) xor (X00 and X40 and X50) xor (X00 and X40 and X52) xor (X00 and X41 and X51) xor (X00 and X41 and X52) xor (X00 and X42 and X51) xor (X0_1 and X40 and X50) xor (X0_1 and X40 and X52) xor (X0_1 and X41 and X50) xor (X0_1 and X42 and X50) xor (X0_1 and X42 and X51) xor (X02 and X40 and X50) xor (X02 and X40 and X51) xor (X02 and X41 and X50) xor (X02 and X41 and X51) xor (X02 and X42 and X50) xor (X02 and X42 and X52) xor (X10 and X40 and X50) xor (X10 and X40 and X52) xor (X10 and X41 and X51) xor (X10 and X41 and X52) xor (X10 and X42 and X51) xor (X11 and X40 and X50) xor (X11 and X40 and X52) xor (X11 and X41 and X50) xor (X11 and X42 and X50) xor (X11 and X42 and X51) xor (X12 and X40 and X50) xor (X12 and X40 and X51) xor (X12 and X41 and X50) xor (X12 and X41 and X51) xor (X12 and X42 and X50) xor (X12 and X42 and X52) xor (X00 and X60) xor (X00 and X61) xor (X02 and X60) xor (X00 and X62) xor (X10 and X60) xor (X10 and X61) xor (X12 and X60) xor (X10 and X62) xor (X00 and X20 and X60) xor (X00 and X20 and X62) xor (X00 and X21 and X61) xor (X00 and X21 and X62) xor (X00 and X22 and X61) xor (X0_1 and X20 and X60) xor (X0_1 and X20 and X62) xor (X0_1 and X21 and X60) xor (X0_1 and X22 and X60) xor (X0_1 and X22 and X61) xor (X02 and X20 and X60) xor (X02 and X20 and X61) xor (X02 and X21 and X60) xor (X02 and X21 and X61) xor (X02 and X22 and X60) xor (X02 and X22 and X62) xor (X30 and X60) xor (X30 and X61) xor (X32 and X60) xor (X30 and X62) xor (X20 and X30 and X60) xor (X20 and X30 and X62) xor (X20 and X31 and X61) xor (X20 and X31 and X62) xor (X20 and X32 and X61) xor (X21 and X30 and X60) xor (X21 and X30 and X62) xor (X21 and X31 and X60) xor (X21 and X32 and X60) xor (X21 and X32 and X61) xor (X22 and X30 and X60) xor (X22 and X30 and X61) xor (X22 and X31 and X60) xor (X22 and X31 and X61) xor (X22 and X32 and X60) xor (X22 and X32 and X62) xor (X00 and X40 and X60) xor (X00 and X40 and X62) xor (X00 and X41 and X61) xor (X00 and X41 and X62) xor (X00 and X42 and X61) xor (X0_1 and X40 and X60) xor (X0_1 and X40 and X62) xor (X0_1 and X41 and X60) xor (X0_1 and X42 and X60) xor (X0_1 and X42 and X61) xor (X02 and X40 and X60) xor (X02 and X40 and X61) xor (X02 and X41 and X60) xor (X02 and X41 and X61) xor (X02 and X42 and X60) xor (X02 and X42 and X62) xor (X10 and X40 and X60) xor (X10 and X40 and X62) xor (X10 and X41 and X61) xor (X10 and X41 and X62) xor (X10 and X42 and X61) xor (X11 and X40 and X60) xor (X11 and X40 and X62) xor (X11 and X41 and X60) xor (X11 and X42 and X60) xor (X11 and X42 and X61) xor (X12 and X40 and X60) xor (X12 and X40 and X61) xor (X12 and X41 and X60) xor (X12 and X41 and X61) xor (X12 and X42 and X60) xor (X12 and X42 and X62) xor (X50 and X60) xor (X50 and X61) xor (X52 and X60) xor (X50 and X62) xor (X00 and X50 and X60) xor (X00 and X50 and X62) xor (X00 and X51 and X61) xor (X00 and X51 and X62) xor (X00 and X52 and X61) xor (X0_1 and X50 and X60) xor (X0_1 and X50 and X62) xor (X0_1 and X51 and X60) xor (X0_1 and X52 and X60) xor (X0_1 and X52 and X61) xor (X02 and X50 and X60) xor (X02 and X50 and X61) xor (X02 and X51 and X60) xor (X02 and X51 and X61) xor (X02 and X52 and X60) xor (X02 and X52 and X62) xor (X40 and X50 and X60) xor (X40 and X50 and X62) xor (X40 and X51 and X61) xor (X40 and X51 and X62) xor (X40 and X52 and X61) xor (X41 and X50 and X60) xor (X41 and X50 and X62) xor (X41 and X51 and X60) xor (X41 and X52 and X60) xor (X41 and X52 and X61) xor (X42 and X50 and X60) xor (X42 and X50 and X61) xor (X42 and X51 and X60) xor (X42 and X51 and X61) xor (X42 and X52 and X60) xor (X42 and X52 and X62) xor (X70) xor (X00 and X70) xor (X00 and X71) xor (X02 and X70) xor (X00 and X72) xor (X10 and X70) xor (X10 and X71) xor (X12 and X70) xor (X10 and X72) xor (X00 and X10 and X70) xor (X00 and X10 and X72) xor (X00 and X11 and X71) xor (X00 and X11 and X72) xor (X00 and X12 and X71) xor (X0_1 and X10 and X70) xor (X0_1 and X10 and X72) xor (X0_1 and X11 and X70) xor (X0_1 and X12 and X70) xor (X0_1 and X12 and X71) xor (X02 and X10 and X70) xor (X02 and X10 and X71) xor (X02 and X11 and X70) xor (X02 and X11 and X71) xor (X02 and X12 and X70) xor (X02 and X12 and X72) xor (X20 and X70) xor (X20 and X71) xor (X22 and X70) xor (X20 and X72) xor (X40 and X70) xor (X40 and X71) xor (X42 and X70) xor (X40 and X72) xor (X00 and X40 and X70) xor (X00 and X40 and X72) xor (X00 and X41 and X71) xor (X00 and X41 and X72) xor (X00 and X42 and X71) xor (X0_1 and X40 and X70) xor (X0_1 and X40 and X72) xor (X0_1 and X41 and X70) xor (X0_1 and X42 and X70) xor (X0_1 and X42 and X71) xor (X02 and X40 and X70) xor (X02 and X40 and X71) xor (X02 and X41 and X70) xor (X02 and X41 and X71) xor (X02 and X42 and X70) xor (X02 and X42 and X72) xor (X50 and X70) xor (X50 and X71) xor (X52 and X70) xor (X50 and X72) xor (X00 and X50 and X70) xor (X00 and X50 and X72) xor (X00 and X51 and X71) xor (X00 and X51 and X72) xor (X00 and X52 and X71) xor (X0_1 and X50 and X70) xor (X0_1 and X50 and X72) xor (X0_1 and X51 and X70) xor (X0_1 and X52 and X70) xor (X0_1 and X52 and X71) xor (X02 and X50 and X70) xor (X02 and X50 and X71) xor (X02 and X51 and X70) xor (X02 and X51 and X71) xor (X02 and X52 and X70) xor (X02 and X52 and X72) xor (X20 and X50 and X70) xor (X20 and X50 and X72) xor (X20 and X51 and X71) xor (X20 and X51 and X72) xor (X20 and X52 and X71) xor (X21 and X50 and X70) xor (X21 and X50 and X72) xor (X21 and X51 and X70) xor (X21 and X52 and X70) xor (X21 and X52 and X71) xor (X22 and X50 and X70) xor (X22 and X50 and X71) xor (X22 and X51 and X70) xor (X22 and X51 and X71) xor (X22 and X52 and X70) xor (X22 and X52 and X72) xor (X40 and X50 and X70) xor (X40 and X50 and X72) xor (X40 and X51 and X71) xor (X40 and X51 and X72) xor (X40 and X52 and X71) xor (X41 and X50 and X70) xor (X41 and X50 and X72) xor (X41 and X51 and X70) xor (X41 and X52 and X70) xor (X41 and X52 and X71) xor (X42 and X50 and X70) xor (X42 and X50 and X71) xor (X42 and X51 and X70) xor (X42 and X51 and X71) xor (X42 and X52 and X70) xor (X42 and X52 and X72) xor (X20 and X60 and X70) xor (X20 and X60 and X72) xor (X20 and X61 and X71) xor (X20 and X61 and X72) xor (X20 and X62 and X71) xor (X21 and X60 and X70) xor (X21 and X60 and X72) xor (X21 and X61 and X70) xor (X21 and X62 and X70) xor (X21 and X62 and X71) xor (X22 and X60 and X70) xor (X22 and X60 and X71) xor (X22 and X61 and X70) xor (X22 and X61 and X71) xor (X22 and X62 and X70) xor (X22 and X62 and X72) xor (X30 and X60 and X70) xor (X30 and X60 and X72) xor (X30 and X61 and X71) xor (X30 and X61 and X72) xor (X30 and X62 and X71) xor (X31 and X60 and X70) xor (X31 and X60 and X72) xor (X31 and X61 and X70) xor (X31 and X62 and X70) xor (X31 and X62 and X71) xor (X32 and X60 and X70) xor (X32 and X60 and X71) xor (X32 and X61 and X70) xor (X32 and X61 and X71) xor (X32 and X62 and X70) xor (X32 and X62 and X72) xor (X40 and X60 and X70) xor (X40 and X60 and X72) xor (X40 and X61 and X71) xor (X40 and X61 and X72) xor (X40 and X62 and X71) xor (X41 and X60 and X70) xor (X41 and X60 and X72) xor (X41 and X61 and X70) xor (X41 and X62 and X70) xor (X41 and X62 and X71) xor (X42 and X60 and X70) xor (X42 and X60 and X71) xor (X42 and X61 and X70) xor (X42 and X61 and X71) xor (X42 and X62 and X70) xor (X42 and X62 and X72));
    F41  <= ((X0_1 and X11) xor (X0_1 and X12) xor (X02 and X11) xor (X0_1 and X13) xor (X21) xor (X31) xor (X0_1 and X31) xor (X0_1 and X32) xor (X02 and X31) xor (X0_1 and X33) xor (X21 and X31) xor (X21 and X32) xor (X22 and X31) xor (X21 and X33) xor (X0_1 and X21 and X31) xor (X0_1 and X21 and X32) xor (X0_1 and X22 and X32) xor (X0_1 and X22 and X33) xor (X0_1 and X23 and X32) xor (X02 and X21 and X32) xor (X02 and X21 and X33) xor (X02 and X22 and X31) xor (X02 and X22 and X33) xor (X02 and X23 and X31) xor (X02 and X23 and X32) xor (X03 and X21 and X32) xor (X03 and X22 and X31) xor (X03 and X22 and X33) xor (X03 and X23 and X31) xor (X03 and X23 and X33) xor (X11 and X21 and X31) xor (X11 and X21 and X32) xor (X11 and X22 and X32) xor (X11 and X22 and X33) xor (X11 and X23 and X32) xor (X12 and X21 and X32) xor (X12 and X21 and X33) xor (X12 and X22 and X31) xor (X12 and X22 and X33) xor (X12 and X23 and X31) xor (X12 and X23 and X32) xor (X13 and X21 and X32) xor (X13 and X22 and X31) xor (X13 and X22 and X33) xor (X13 and X23 and X31) xor (X13 and X23 and X33) xor (X11 and X41) xor (X11 and X42) xor (X12 and X41) xor (X11 and X43) xor (X0_1 and X11 and X41) xor (X0_1 and X11 and X42) xor (X0_1 and X12 and X42) xor (X0_1 and X12 and X43) xor (X0_1 and X13 and X42) xor (X02 and X11 and X42) xor (X02 and X11 and X43) xor (X02 and X12 and X41) xor (X02 and X12 and X43) xor (X02 and X13 and X41) xor (X02 and X13 and X42) xor (X03 and X11 and X42) xor (X03 and X12 and X41) xor (X03 and X12 and X43) xor (X03 and X13 and X41) xor (X03 and X13 and X43) xor (X31 and X41) xor (X31 and X42) xor (X32 and X41) xor (X31 and X43) xor (X0_1 and X31 and X41) xor (X0_1 and X31 and X42) xor (X0_1 and X32 and X42) xor (X0_1 and X32 and X43) xor (X0_1 and X33 and X42) xor (X02 and X31 and X42) xor (X02 and X31 and X43) xor (X02 and X32 and X41) xor (X02 and X32 and X43) xor (X02 and X33 and X41) xor (X02 and X33 and X42) xor (X03 and X31 and X42) xor (X03 and X32 and X41) xor (X03 and X32 and X43) xor (X03 and X33 and X41) xor (X03 and X33 and X43) xor (X11 and X31 and X41) xor (X11 and X31 and X42) xor (X11 and X32 and X42) xor (X11 and X32 and X43) xor (X11 and X33 and X42) xor (X12 and X31 and X42) xor (X12 and X31 and X43) xor (X12 and X32 and X41) xor (X12 and X32 and X43) xor (X12 and X33 and X41) xor (X12 and X33 and X42) xor (X13 and X31 and X42) xor (X13 and X32 and X41) xor (X13 and X32 and X43) xor (X13 and X33 and X41) xor (X13 and X33 and X43) xor (X21 and X31 and X41) xor (X21 and X31 and X42) xor (X21 and X32 and X42) xor (X21 and X32 and X43) xor (X21 and X33 and X42) xor (X22 and X31 and X42) xor (X22 and X31 and X43) xor (X22 and X32 and X41) xor (X22 and X32 and X43) xor (X22 and X33 and X41) xor (X22 and X33 and X42) xor (X23 and X31 and X42) xor (X23 and X32 and X41) xor (X23 and X32 and X43) xor (X23 and X33 and X41) xor (X23 and X33 and X43) xor (X51) xor (X11 and X51) xor (X11 and X52) xor (X12 and X51) xor (X11 and X53) xor (X0_1 and X11 and X51) xor (X0_1 and X11 and X52) xor (X0_1 and X12 and X52) xor (X0_1 and X12 and X53) xor (X0_1 and X13 and X52) xor (X02 and X11 and X52) xor (X02 and X11 and X53) xor (X02 and X12 and X51) xor (X02 and X12 and X53) xor (X02 and X13 and X51) xor (X02 and X13 and X52) xor (X03 and X11 and X52) xor (X03 and X12 and X51) xor (X03 and X12 and X53) xor (X03 and X13 and X51) xor (X03 and X13 and X53) xor (X0_1 and X21 and X51) xor (X0_1 and X21 and X52) xor (X0_1 and X22 and X52) xor (X0_1 and X22 and X53) xor (X0_1 and X23 and X52) xor (X02 and X21 and X52) xor (X02 and X21 and X53) xor (X02 and X22 and X51) xor (X02 and X22 and X53) xor (X02 and X23 and X51) xor (X02 and X23 and X52) xor (X03 and X21 and X52) xor (X03 and X22 and X51) xor (X03 and X22 and X53) xor (X03 and X23 and X51) xor (X03 and X23 and X53) xor (X11 and X21 and X51) xor (X11 and X21 and X52) xor (X11 and X22 and X52) xor (X11 and X22 and X53) xor (X11 and X23 and X52) xor (X12 and X21 and X52) xor (X12 and X21 and X53) xor (X12 and X22 and X51) xor (X12 and X22 and X53) xor (X12 and X23 and X51) xor (X12 and X23 and X52) xor (X13 and X21 and X52) xor (X13 and X22 and X51) xor (X13 and X22 and X53) xor (X13 and X23 and X51) xor (X13 and X23 and X53) xor (X31 and X51) xor (X31 and X52) xor (X32 and X51) xor (X31 and X53) xor (X11 and X31 and X51) xor (X11 and X31 and X52) xor (X11 and X32 and X52) xor (X11 and X32 and X53) xor (X11 and X33 and X52) xor (X12 and X31 and X52) xor (X12 and X31 and X53) xor (X12 and X32 and X51) xor (X12 and X32 and X53) xor (X12 and X33 and X51) xor (X12 and X33 and X52) xor (X13 and X31 and X52) xor (X13 and X32 and X51) xor (X13 and X32 and X53) xor (X13 and X33 and X51) xor (X13 and X33 and X53) xor (X21 and X31 and X51) xor (X21 and X31 and X52) xor (X21 and X32 and X52) xor (X21 and X32 and X53) xor (X21 and X33 and X52) xor (X22 and X31 and X52) xor (X22 and X31 and X53) xor (X22 and X32 and X51) xor (X22 and X32 and X53) xor (X22 and X33 and X51) xor (X22 and X33 and X52) xor (X23 and X31 and X52) xor (X23 and X32 and X51) xor (X23 and X32 and X53) xor (X23 and X33 and X51) xor (X23 and X33 and X53) xor (X41 and X51) xor (X41 and X52) xor (X42 and X51) xor (X41 and X53) xor (X0_1 and X41 and X51) xor (X0_1 and X41 and X52) xor (X0_1 and X42 and X52) xor (X0_1 and X42 and X53) xor (X0_1 and X43 and X52) xor (X02 and X41 and X52) xor (X02 and X41 and X53) xor (X02 and X42 and X51) xor (X02 and X42 and X53) xor (X02 and X43 and X51) xor (X02 and X43 and X52) xor (X03 and X41 and X52) xor (X03 and X42 and X51) xor (X03 and X42 and X53) xor (X03 and X43 and X51) xor (X03 and X43 and X53) xor (X11 and X41 and X51) xor (X11 and X41 and X52) xor (X11 and X42 and X52) xor (X11 and X42 and X53) xor (X11 and X43 and X52) xor (X12 and X41 and X52) xor (X12 and X41 and X53) xor (X12 and X42 and X51) xor (X12 and X42 and X53) xor (X12 and X43 and X51) xor (X12 and X43 and X52) xor (X13 and X41 and X52) xor (X13 and X42 and X51) xor (X13 and X42 and X53) xor (X13 and X43 and X51) xor (X13 and X43 and X53) xor (X0_1 and X61) xor (X0_1 and X62) xor (X02 and X61) xor (X0_1 and X63) xor (X11 and X61) xor (X11 and X62) xor (X12 and X61) xor (X11 and X63) xor (X0_1 and X21 and X61) xor (X0_1 and X21 and X62) xor (X0_1 and X22 and X62) xor (X0_1 and X22 and X63) xor (X0_1 and X23 and X62) xor (X02 and X21 and X62) xor (X02 and X21 and X63) xor (X02 and X22 and X61) xor (X02 and X22 and X63) xor (X02 and X23 and X61) xor (X02 and X23 and X62) xor (X03 and X21 and X62) xor (X03 and X22 and X61) xor (X03 and X22 and X63) xor (X03 and X23 and X61) xor (X03 and X23 and X63) xor (X31 and X61) xor (X31 and X62) xor (X32 and X61) xor (X31 and X63) xor (X21 and X31 and X61) xor (X21 and X31 and X62) xor (X21 and X32 and X62) xor (X21 and X32 and X63) xor (X21 and X33 and X62) xor (X22 and X31 and X62) xor (X22 and X31 and X63) xor (X22 and X32 and X61) xor (X22 and X32 and X63) xor (X22 and X33 and X61) xor (X22 and X33 and X62) xor (X23 and X31 and X62) xor (X23 and X32 and X61) xor (X23 and X32 and X63) xor (X23 and X33 and X61) xor (X23 and X33 and X63) xor (X0_1 and X41 and X61) xor (X0_1 and X41 and X62) xor (X0_1 and X42 and X62) xor (X0_1 and X42 and X63) xor (X0_1 and X43 and X62) xor (X02 and X41 and X62) xor (X02 and X41 and X63) xor (X02 and X42 and X61) xor (X02 and X42 and X63) xor (X02 and X43 and X61) xor (X02 and X43 and X62) xor (X03 and X41 and X62) xor (X03 and X42 and X61) xor (X03 and X42 and X63) xor (X03 and X43 and X61) xor (X03 and X43 and X63) xor (X11 and X41 and X61) xor (X11 and X41 and X62) xor (X11 and X42 and X62) xor (X11 and X42 and X63) xor (X11 and X43 and X62) xor (X12 and X41 and X62) xor (X12 and X41 and X63) xor (X12 and X42 and X61) xor (X12 and X42 and X63) xor (X12 and X43 and X61) xor (X12 and X43 and X62) xor (X13 and X41 and X62) xor (X13 and X42 and X61) xor (X13 and X42 and X63) xor (X13 and X43 and X61) xor (X13 and X43 and X63) xor (X51 and X61) xor (X51 and X62) xor (X52 and X61) xor (X51 and X63) xor (X0_1 and X51 and X61) xor (X0_1 and X51 and X62) xor (X0_1 and X52 and X62) xor (X0_1 and X52 and X63) xor (X0_1 and X53 and X62) xor (X02 and X51 and X62) xor (X02 and X51 and X63) xor (X02 and X52 and X61) xor (X02 and X52 and X63) xor (X02 and X53 and X61) xor (X02 and X53 and X62) xor (X03 and X51 and X62) xor (X03 and X52 and X61) xor (X03 and X52 and X63) xor (X03 and X53 and X61) xor (X03 and X53 and X63) xor (X41 and X51 and X61) xor (X41 and X51 and X62) xor (X41 and X52 and X62) xor (X41 and X52 and X63) xor (X41 and X53 and X62) xor (X42 and X51 and X62) xor (X42 and X51 and X63) xor (X42 and X52 and X61) xor (X42 and X52 and X63) xor (X42 and X53 and X61) xor (X42 and X53 and X62) xor (X43 and X51 and X62) xor (X43 and X52 and X61) xor (X43 and X52 and X63) xor (X43 and X53 and X61) xor (X43 and X53 and X63) xor (X71) xor (X0_1 and X71) xor (X0_1 and X72) xor (X02 and X71) xor (X0_1 and X73) xor (X11 and X71) xor (X11 and X72) xor (X12 and X71) xor (X11 and X73) xor (X0_1 and X11 and X71) xor (X0_1 and X11 and X72) xor (X0_1 and X12 and X72) xor (X0_1 and X12 and X73) xor (X0_1 and X13 and X72) xor (X02 and X11 and X72) xor (X02 and X11 and X73) xor (X02 and X12 and X71) xor (X02 and X12 and X73) xor (X02 and X13 and X71) xor (X02 and X13 and X72) xor (X03 and X11 and X72) xor (X03 and X12 and X71) xor (X03 and X12 and X73) xor (X03 and X13 and X71) xor (X03 and X13 and X73) xor (X21 and X71) xor (X21 and X72) xor (X22 and X71) xor (X21 and X73) xor (X41 and X71) xor (X41 and X72) xor (X42 and X71) xor (X41 and X73) xor (X0_1 and X41 and X71) xor (X0_1 and X41 and X72) xor (X0_1 and X42 and X72) xor (X0_1 and X42 and X73) xor (X0_1 and X43 and X72) xor (X02 and X41 and X72) xor (X02 and X41 and X73) xor (X02 and X42 and X71) xor (X02 and X42 and X73) xor (X02 and X43 and X71) xor (X02 and X43 and X72) xor (X03 and X41 and X72) xor (X03 and X42 and X71) xor (X03 and X42 and X73) xor (X03 and X43 and X71) xor (X03 and X43 and X73) xor (X51 and X71) xor (X51 and X72) xor (X52 and X71) xor (X51 and X73) xor (X0_1 and X51 and X71) xor (X0_1 and X51 and X72) xor (X0_1 and X52 and X72) xor (X0_1 and X52 and X73) xor (X0_1 and X53 and X72) xor (X02 and X51 and X72) xor (X02 and X51 and X73) xor (X02 and X52 and X71) xor (X02 and X52 and X73) xor (X02 and X53 and X71) xor (X02 and X53 and X72) xor (X03 and X51 and X72) xor (X03 and X52 and X71) xor (X03 and X52 and X73) xor (X03 and X53 and X71) xor (X03 and X53 and X73) xor (X21 and X51 and X71) xor (X21 and X51 and X72) xor (X21 and X52 and X72) xor (X21 and X52 and X73) xor (X21 and X53 and X72) xor (X22 and X51 and X72) xor (X22 and X51 and X73) xor (X22 and X52 and X71) xor (X22 and X52 and X73) xor (X22 and X53 and X71) xor (X22 and X53 and X72) xor (X23 and X51 and X72) xor (X23 and X52 and X71) xor (X23 and X52 and X73) xor (X23 and X53 and X71) xor (X23 and X53 and X73) xor (X41 and X51 and X71) xor (X41 and X51 and X72) xor (X41 and X52 and X72) xor (X41 and X52 and X73) xor (X41 and X53 and X72) xor (X42 and X51 and X72) xor (X42 and X51 and X73) xor (X42 and X52 and X71) xor (X42 and X52 and X73) xor (X42 and X53 and X71) xor (X42 and X53 and X72) xor (X43 and X51 and X72) xor (X43 and X52 and X71) xor (X43 and X52 and X73) xor (X43 and X53 and X71) xor (X43 and X53 and X73) xor (X21 and X61 and X71) xor (X21 and X61 and X72) xor (X21 and X62 and X72) xor (X21 and X62 and X73) xor (X21 and X63 and X72) xor (X22 and X61 and X72) xor (X22 and X61 and X73) xor (X22 and X62 and X71) xor (X22 and X62 and X73) xor (X22 and X63 and X71) xor (X22 and X63 and X72) xor (X23 and X61 and X72) xor (X23 and X62 and X71) xor (X23 and X62 and X73) xor (X23 and X63 and X71) xor (X23 and X63 and X73) xor (X31 and X61 and X71) xor (X31 and X61 and X72) xor (X31 and X62 and X72) xor (X31 and X62 and X73) xor (X31 and X63 and X72) xor (X32 and X61 and X72) xor (X32 and X61 and X73) xor (X32 and X62 and X71) xor (X32 and X62 and X73) xor (X32 and X63 and X71) xor (X32 and X63 and X72) xor (X33 and X61 and X72) xor (X33 and X62 and X71) xor (X33 and X62 and X73) xor (X33 and X63 and X71) xor (X33 and X63 and X73) xor (X41 and X61 and X71) xor (X41 and X61 and X72) xor (X41 and X62 and X72) xor (X41 and X62 and X73) xor (X41 and X63 and X72) xor (X42 and X61 and X72) xor (X42 and X61 and X73) xor (X42 and X62 and X71) xor (X42 and X62 and X73) xor (X42 and X63 and X71) xor (X42 and X63 and X72) xor (X43 and X61 and X72) xor (X43 and X62 and X71) xor (X43 and X62 and X73) xor (X43 and X63 and X71) xor (X43 and X63 and X73));
    F42  <= ((X02 and X12) xor (X00 and X13) xor (X02 and X13) xor (X03 and X12) xor (X22) xor (X32) xor (X02 and X32) xor (X00 and X33) xor (X02 and X33) xor (X03 and X32) xor (X22 and X32) xor (X20 and X33) xor (X22 and X33) xor (X23 and X32) xor (X00 and X20 and X33) xor (X00 and X22 and X30) xor (X00 and X22 and X32) xor (X00 and X22 and X33) xor (X00 and X23 and X30) xor (X00 and X23 and X32) xor (X02 and X20 and X32) xor (X02 and X20 and X33) xor (X02 and X23 and X30) xor (X02 and X23 and X33) xor (X03 and X20 and X30) xor (X03 and X20 and X32) xor (X03 and X20 and X33) xor (X03 and X22 and X30) xor (X03 and X22 and X32) xor (X03 and X23 and X32) xor (X10 and X20 and X33) xor (X10 and X22 and X30) xor (X10 and X22 and X32) xor (X10 and X22 and X33) xor (X10 and X23 and X30) xor (X10 and X23 and X32) xor (X12 and X20 and X32) xor (X12 and X20 and X33) xor (X12 and X23 and X30) xor (X12 and X23 and X33) xor (X13 and X20 and X30) xor (X13 and X20 and X32) xor (X13 and X20 and X33) xor (X13 and X22 and X30) xor (X13 and X22 and X32) xor (X13 and X23 and X32) xor (X12 and X42) xor (X10 and X43) xor (X12 and X43) xor (X13 and X42) xor (X00 and X10 and X43) xor (X00 and X12 and X40) xor (X00 and X12 and X42) xor (X00 and X12 and X43) xor (X00 and X13 and X40) xor (X00 and X13 and X42) xor (X02 and X10 and X42) xor (X02 and X10 and X43) xor (X02 and X13 and X40) xor (X02 and X13 and X43) xor (X03 and X10 and X40) xor (X03 and X10 and X42) xor (X03 and X10 and X43) xor (X03 and X12 and X40) xor (X03 and X12 and X42) xor (X03 and X13 and X42) xor (X32 and X42) xor (X30 and X43) xor (X32 and X43) xor (X33 and X42) xor (X00 and X30 and X43) xor (X00 and X32 and X40) xor (X00 and X32 and X42) xor (X00 and X32 and X43) xor (X00 and X33 and X40) xor (X00 and X33 and X42) xor (X02 and X30 and X42) xor (X02 and X30 and X43) xor (X02 and X33 and X40) xor (X02 and X33 and X43) xor (X03 and X30 and X40) xor (X03 and X30 and X42) xor (X03 and X30 and X43) xor (X03 and X32 and X40) xor (X03 and X32 and X42) xor (X03 and X33 and X42) xor (X10 and X30 and X43) xor (X10 and X32 and X40) xor (X10 and X32 and X42) xor (X10 and X32 and X43) xor (X10 and X33 and X40) xor (X10 and X33 and X42) xor (X12 and X30 and X42) xor (X12 and X30 and X43) xor (X12 and X33 and X40) xor (X12 and X33 and X43) xor (X13 and X30 and X40) xor (X13 and X30 and X42) xor (X13 and X30 and X43) xor (X13 and X32 and X40) xor (X13 and X32 and X42) xor (X13 and X33 and X42) xor (X20 and X30 and X43) xor (X20 and X32 and X40) xor (X20 and X32 and X42) xor (X20 and X32 and X43) xor (X20 and X33 and X40) xor (X20 and X33 and X42) xor (X22 and X30 and X42) xor (X22 and X30 and X43) xor (X22 and X33 and X40) xor (X22 and X33 and X43) xor (X23 and X30 and X40) xor (X23 and X30 and X42) xor (X23 and X30 and X43) xor (X23 and X32 and X40) xor (X23 and X32 and X42) xor (X23 and X33 and X42) xor (X52) xor (X12 and X52) xor (X10 and X53) xor (X12 and X53) xor (X13 and X52) xor (X00 and X10 and X53) xor (X00 and X12 and X50) xor (X00 and X12 and X52) xor (X00 and X12 and X53) xor (X00 and X13 and X50) xor (X00 and X13 and X52) xor (X02 and X10 and X52) xor (X02 and X10 and X53) xor (X02 and X13 and X50) xor (X02 and X13 and X53) xor (X03 and X10 and X50) xor (X03 and X10 and X52) xor (X03 and X10 and X53) xor (X03 and X12 and X50) xor (X03 and X12 and X52) xor (X03 and X13 and X52) xor (X00 and X20 and X53) xor (X00 and X22 and X50) xor (X00 and X22 and X52) xor (X00 and X22 and X53) xor (X00 and X23 and X50) xor (X00 and X23 and X52) xor (X02 and X20 and X52) xor (X02 and X20 and X53) xor (X02 and X23 and X50) xor (X02 and X23 and X53) xor (X03 and X20 and X50) xor (X03 and X20 and X52) xor (X03 and X20 and X53) xor (X03 and X22 and X50) xor (X03 and X22 and X52) xor (X03 and X23 and X52) xor (X10 and X20 and X53) xor (X10 and X22 and X50) xor (X10 and X22 and X52) xor (X10 and X22 and X53) xor (X10 and X23 and X50) xor (X10 and X23 and X52) xor (X12 and X20 and X52) xor (X12 and X20 and X53) xor (X12 and X23 and X50) xor (X12 and X23 and X53) xor (X13 and X20 and X50) xor (X13 and X20 and X52) xor (X13 and X20 and X53) xor (X13 and X22 and X50) xor (X13 and X22 and X52) xor (X13 and X23 and X52) xor (X32 and X52) xor (X30 and X53) xor (X32 and X53) xor (X33 and X52) xor (X10 and X30 and X53) xor (X10 and X32 and X50) xor (X10 and X32 and X52) xor (X10 and X32 and X53) xor (X10 and X33 and X50) xor (X10 and X33 and X52) xor (X12 and X30 and X52) xor (X12 and X30 and X53) xor (X12 and X33 and X50) xor (X12 and X33 and X53) xor (X13 and X30 and X50) xor (X13 and X30 and X52) xor (X13 and X30 and X53) xor (X13 and X32 and X50) xor (X13 and X32 and X52) xor (X13 and X33 and X52) xor (X20 and X30 and X53) xor (X20 and X32 and X50) xor (X20 and X32 and X52) xor (X20 and X32 and X53) xor (X20 and X33 and X50) xor (X20 and X33 and X52) xor (X22 and X30 and X52) xor (X22 and X30 and X53) xor (X22 and X33 and X50) xor (X22 and X33 and X53) xor (X23 and X30 and X50) xor (X23 and X30 and X52) xor (X23 and X30 and X53) xor (X23 and X32 and X50) xor (X23 and X32 and X52) xor (X23 and X33 and X52) xor (X42 and X52) xor (X40 and X53) xor (X42 and X53) xor (X43 and X52) xor (X00 and X40 and X53) xor (X00 and X42 and X50) xor (X00 and X42 and X52) xor (X00 and X42 and X53) xor (X00 and X43 and X50) xor (X00 and X43 and X52) xor (X02 and X40 and X52) xor (X02 and X40 and X53) xor (X02 and X43 and X50) xor (X02 and X43 and X53) xor (X03 and X40 and X50) xor (X03 and X40 and X52) xor (X03 and X40 and X53) xor (X03 and X42 and X50) xor (X03 and X42 and X52) xor (X03 and X43 and X52) xor (X10 and X40 and X53) xor (X10 and X42 and X50) xor (X10 and X42 and X52) xor (X10 and X42 and X53) xor (X10 and X43 and X50) xor (X10 and X43 and X52) xor (X12 and X40 and X52) xor (X12 and X40 and X53) xor (X12 and X43 and X50) xor (X12 and X43 and X53) xor (X13 and X40 and X50) xor (X13 and X40 and X52) xor (X13 and X40 and X53) xor (X13 and X42 and X50) xor (X13 and X42 and X52) xor (X13 and X43 and X52) xor (X02 and X62) xor (X00 and X63) xor (X02 and X63) xor (X03 and X62) xor (X12 and X62) xor (X10 and X63) xor (X12 and X63) xor (X13 and X62) xor (X00 and X20 and X63) xor (X00 and X22 and X60) xor (X00 and X22 and X62) xor (X00 and X22 and X63) xor (X00 and X23 and X60) xor (X00 and X23 and X62) xor (X02 and X20 and X62) xor (X02 and X20 and X63) xor (X02 and X23 and X60) xor (X02 and X23 and X63) xor (X03 and X20 and X60) xor (X03 and X20 and X62) xor (X03 and X20 and X63) xor (X03 and X22 and X60) xor (X03 and X22 and X62) xor (X03 and X23 and X62) xor (X32 and X62) xor (X30 and X63) xor (X32 and X63) xor (X33 and X62) xor (X20 and X30 and X63) xor (X20 and X32 and X60) xor (X20 and X32 and X62) xor (X20 and X32 and X63) xor (X20 and X33 and X60) xor (X20 and X33 and X62) xor (X22 and X30 and X62) xor (X22 and X30 and X63) xor (X22 and X33 and X60) xor (X22 and X33 and X63) xor (X23 and X30 and X60) xor (X23 and X30 and X62) xor (X23 and X30 and X63) xor (X23 and X32 and X60) xor (X23 and X32 and X62) xor (X23 and X33 and X62) xor (X00 and X40 and X63) xor (X00 and X42 and X60) xor (X00 and X42 and X62) xor (X00 and X42 and X63) xor (X00 and X43 and X60) xor (X00 and X43 and X62) xor (X02 and X40 and X62) xor (X02 and X40 and X63) xor (X02 and X43 and X60) xor (X02 and X43 and X63) xor (X03 and X40 and X60) xor (X03 and X40 and X62) xor (X03 and X40 and X63) xor (X03 and X42 and X60) xor (X03 and X42 and X62) xor (X03 and X43 and X62) xor (X10 and X40 and X63) xor (X10 and X42 and X60) xor (X10 and X42 and X62) xor (X10 and X42 and X63) xor (X10 and X43 and X60) xor (X10 and X43 and X62) xor (X12 and X40 and X62) xor (X12 and X40 and X63) xor (X12 and X43 and X60) xor (X12 and X43 and X63) xor (X13 and X40 and X60) xor (X13 and X40 and X62) xor (X13 and X40 and X63) xor (X13 and X42 and X60) xor (X13 and X42 and X62) xor (X13 and X43 and X62) xor (X52 and X62) xor (X50 and X63) xor (X52 and X63) xor (X53 and X62) xor (X00 and X50 and X63) xor (X00 and X52 and X60) xor (X00 and X52 and X62) xor (X00 and X52 and X63) xor (X00 and X53 and X60) xor (X00 and X53 and X62) xor (X02 and X50 and X62) xor (X02 and X50 and X63) xor (X02 and X53 and X60) xor (X02 and X53 and X63) xor (X03 and X50 and X60) xor (X03 and X50 and X62) xor (X03 and X50 and X63) xor (X03 and X52 and X60) xor (X03 and X52 and X62) xor (X03 and X53 and X62) xor (X40 and X50 and X63) xor (X40 and X52 and X60) xor (X40 and X52 and X62) xor (X40 and X52 and X63) xor (X40 and X53 and X60) xor (X40 and X53 and X62) xor (X42 and X50 and X62) xor (X42 and X50 and X63) xor (X42 and X53 and X60) xor (X42 and X53 and X63) xor (X43 and X50 and X60) xor (X43 and X50 and X62) xor (X43 and X50 and X63) xor (X43 and X52 and X60) xor (X43 and X52 and X62) xor (X43 and X53 and X62) xor (X72) xor (X02 and X72) xor (X00 and X73) xor (X02 and X73) xor (X03 and X72) xor (X12 and X72) xor (X10 and X73) xor (X12 and X73) xor (X13 and X72) xor (X00 and X10 and X73) xor (X00 and X12 and X70) xor (X00 and X12 and X72) xor (X00 and X12 and X73) xor (X00 and X13 and X70) xor (X00 and X13 and X72) xor (X02 and X10 and X72) xor (X02 and X10 and X73) xor (X02 and X13 and X70) xor (X02 and X13 and X73) xor (X03 and X10 and X70) xor (X03 and X10 and X72) xor (X03 and X10 and X73) xor (X03 and X12 and X70) xor (X03 and X12 and X72) xor (X03 and X13 and X72) xor (X22 and X72) xor (X20 and X73) xor (X22 and X73) xor (X23 and X72) xor (X42 and X72) xor (X40 and X73) xor (X42 and X73) xor (X43 and X72) xor (X00 and X40 and X73) xor (X00 and X42 and X70) xor (X00 and X42 and X72) xor (X00 and X42 and X73) xor (X00 and X43 and X70) xor (X00 and X43 and X72) xor (X02 and X40 and X72) xor (X02 and X40 and X73) xor (X02 and X43 and X70) xor (X02 and X43 and X73) xor (X03 and X40 and X70) xor (X03 and X40 and X72) xor (X03 and X40 and X73) xor (X03 and X42 and X70) xor (X03 and X42 and X72) xor (X03 and X43 and X72) xor (X52 and X72) xor (X50 and X73) xor (X52 and X73) xor (X53 and X72) xor (X00 and X50 and X73) xor (X00 and X52 and X70) xor (X00 and X52 and X72) xor (X00 and X52 and X73) xor (X00 and X53 and X70) xor (X00 and X53 and X72) xor (X02 and X50 and X72) xor (X02 and X50 and X73) xor (X02 and X53 and X70) xor (X02 and X53 and X73) xor (X03 and X50 and X70) xor (X03 and X50 and X72) xor (X03 and X50 and X73) xor (X03 and X52 and X70) xor (X03 and X52 and X72) xor (X03 and X53 and X72) xor (X20 and X50 and X73) xor (X20 and X52 and X70) xor (X20 and X52 and X72) xor (X20 and X52 and X73) xor (X20 and X53 and X70) xor (X20 and X53 and X72) xor (X22 and X50 and X72) xor (X22 and X50 and X73) xor (X22 and X53 and X70) xor (X22 and X53 and X73) xor (X23 and X50 and X70) xor (X23 and X50 and X72) xor (X23 and X50 and X73) xor (X23 and X52 and X70) xor (X23 and X52 and X72) xor (X23 and X53 and X72) xor (X40 and X50 and X73) xor (X40 and X52 and X70) xor (X40 and X52 and X72) xor (X40 and X52 and X73) xor (X40 and X53 and X70) xor (X40 and X53 and X72) xor (X42 and X50 and X72) xor (X42 and X50 and X73) xor (X42 and X53 and X70) xor (X42 and X53 and X73) xor (X43 and X50 and X70) xor (X43 and X50 and X72) xor (X43 and X50 and X73) xor (X43 and X52 and X70) xor (X43 and X52 and X72) xor (X43 and X53 and X72) xor (X20 and X60 and X73) xor (X20 and X62 and X70) xor (X20 and X62 and X72) xor (X20 and X62 and X73) xor (X20 and X63 and X70) xor (X20 and X63 and X72) xor (X22 and X60 and X72) xor (X22 and X60 and X73) xor (X22 and X63 and X70) xor (X22 and X63 and X73) xor (X23 and X60 and X70) xor (X23 and X60 and X72) xor (X23 and X60 and X73) xor (X23 and X62 and X70) xor (X23 and X62 and X72) xor (X23 and X63 and X72) xor (X30 and X60 and X73) xor (X30 and X62 and X70) xor (X30 and X62 and X72) xor (X30 and X62 and X73) xor (X30 and X63 and X70) xor (X30 and X63 and X72) xor (X32 and X60 and X72) xor (X32 and X60 and X73) xor (X32 and X63 and X70) xor (X32 and X63 and X73) xor (X33 and X60 and X70) xor (X33 and X60 and X72) xor (X33 and X60 and X73) xor (X33 and X62 and X70) xor (X33 and X62 and X72) xor (X33 and X63 and X72) xor (X40 and X60 and X73) xor (X40 and X62 and X70) xor (X40 and X62 and X72) xor (X40 and X62 and X73) xor (X40 and X63 and X70) xor (X40 and X63 and X72) xor (X42 and X60 and X72) xor (X42 and X60 and X73) xor (X42 and X63 and X70) xor (X42 and X63 and X73) xor (X43 and X60 and X70) xor (X43 and X60 and X72) xor (X43 and X60 and X73) xor (X43 and X62 and X70) xor (X43 and X62 and X72) xor (X43 and X63 and X72));
    F43  <= ((X03 and X13) xor (X03 and X10) xor (X03 and X11) xor (X0_1 and X10) xor (X23) xor (X33) xor (X03 and X33) xor (X03 and X30) xor (X03 and X31) xor (X0_1 and X30) xor (X23 and X33) xor (X23 and X30) xor (X23 and X31) xor (X21 and X30) xor (X00 and X20 and X31) xor (X00 and X21 and X30) xor (X00 and X21 and X33) xor (X00 and X23 and X31) xor (X00 and X23 and X33) xor (X0_1 and X20 and X31) xor (X0_1 and X20 and X33) xor (X0_1 and X21 and X33) xor (X0_1 and X23 and X30) xor (X0_1 and X23 and X31) xor (X0_1 and X23 and X33) xor (X03 and X20 and X31) xor (X03 and X21 and X30) xor (X03 and X21 and X31) xor (X03 and X21 and X33) xor (X03 and X23 and X30) xor (X10 and X20 and X31) xor (X10 and X21 and X30) xor (X10 and X21 and X33) xor (X10 and X23 and X31) xor (X10 and X23 and X33) xor (X11 and X20 and X31) xor (X11 and X20 and X33) xor (X11 and X21 and X33) xor (X11 and X23 and X30) xor (X11 and X23 and X31) xor (X11 and X23 and X33) xor (X13 and X20 and X31) xor (X13 and X21 and X30) xor (X13 and X21 and X31) xor (X13 and X21 and X33) xor (X13 and X23 and X30) xor (X13 and X43) xor (X13 and X40) xor (X13 and X41) xor (X11 and X40) xor (X00 and X10 and X41) xor (X00 and X11 and X40) xor (X00 and X11 and X43) xor (X00 and X13 and X41) xor (X00 and X13 and X43) xor (X0_1 and X10 and X41) xor (X0_1 and X10 and X43) xor (X0_1 and X11 and X43) xor (X0_1 and X13 and X40) xor (X0_1 and X13 and X41) xor (X0_1 and X13 and X43) xor (X03 and X10 and X41) xor (X03 and X11 and X40) xor (X03 and X11 and X41) xor (X03 and X11 and X43) xor (X03 and X13 and X40) xor (X33 and X43) xor (X33 and X40) xor (X33 and X41) xor (X31 and X40) xor (X00 and X30 and X41) xor (X00 and X31 and X40) xor (X00 and X31 and X43) xor (X00 and X33 and X41) xor (X00 and X33 and X43) xor (X0_1 and X30 and X41) xor (X0_1 and X30 and X43) xor (X0_1 and X31 and X43) xor (X0_1 and X33 and X40) xor (X0_1 and X33 and X41) xor (X0_1 and X33 and X43) xor (X03 and X30 and X41) xor (X03 and X31 and X40) xor (X03 and X31 and X41) xor (X03 and X31 and X43) xor (X03 and X33 and X40) xor (X10 and X30 and X41) xor (X10 and X31 and X40) xor (X10 and X31 and X43) xor (X10 and X33 and X41) xor (X10 and X33 and X43) xor (X11 and X30 and X41) xor (X11 and X30 and X43) xor (X11 and X31 and X43) xor (X11 and X33 and X40) xor (X11 and X33 and X41) xor (X11 and X33 and X43) xor (X13 and X30 and X41) xor (X13 and X31 and X40) xor (X13 and X31 and X41) xor (X13 and X31 and X43) xor (X13 and X33 and X40) xor (X20 and X30 and X41) xor (X20 and X31 and X40) xor (X20 and X31 and X43) xor (X20 and X33 and X41) xor (X20 and X33 and X43) xor (X21 and X30 and X41) xor (X21 and X30 and X43) xor (X21 and X31 and X43) xor (X21 and X33 and X40) xor (X21 and X33 and X41) xor (X21 and X33 and X43) xor (X23 and X30 and X41) xor (X23 and X31 and X40) xor (X23 and X31 and X41) xor (X23 and X31 and X43) xor (X23 and X33 and X40) xor (X53) xor (X13 and X53) xor (X13 and X50) xor (X13 and X51) xor (X11 and X50) xor (X00 and X10 and X51) xor (X00 and X11 and X50) xor (X00 and X11 and X53) xor (X00 and X13 and X51) xor (X00 and X13 and X53) xor (X0_1 and X10 and X51) xor (X0_1 and X10 and X53) xor (X0_1 and X11 and X53) xor (X0_1 and X13 and X50) xor (X0_1 and X13 and X51) xor (X0_1 and X13 and X53) xor (X03 and X10 and X51) xor (X03 and X11 and X50) xor (X03 and X11 and X51) xor (X03 and X11 and X53) xor (X03 and X13 and X50) xor (X00 and X20 and X51) xor (X00 and X21 and X50) xor (X00 and X21 and X53) xor (X00 and X23 and X51) xor (X00 and X23 and X53) xor (X0_1 and X20 and X51) xor (X0_1 and X20 and X53) xor (X0_1 and X21 and X53) xor (X0_1 and X23 and X50) xor (X0_1 and X23 and X51) xor (X0_1 and X23 and X53) xor (X03 and X20 and X51) xor (X03 and X21 and X50) xor (X03 and X21 and X51) xor (X03 and X21 and X53) xor (X03 and X23 and X50) xor (X10 and X20 and X51) xor (X10 and X21 and X50) xor (X10 and X21 and X53) xor (X10 and X23 and X51) xor (X10 and X23 and X53) xor (X11 and X20 and X51) xor (X11 and X20 and X53) xor (X11 and X21 and X53) xor (X11 and X23 and X50) xor (X11 and X23 and X51) xor (X11 and X23 and X53) xor (X13 and X20 and X51) xor (X13 and X21 and X50) xor (X13 and X21 and X51) xor (X13 and X21 and X53) xor (X13 and X23 and X50) xor (X33 and X53) xor (X33 and X50) xor (X33 and X51) xor (X31 and X50) xor (X10 and X30 and X51) xor (X10 and X31 and X50) xor (X10 and X31 and X53) xor (X10 and X33 and X51) xor (X10 and X33 and X53) xor (X11 and X30 and X51) xor (X11 and X30 and X53) xor (X11 and X31 and X53) xor (X11 and X33 and X50) xor (X11 and X33 and X51) xor (X11 and X33 and X53) xor (X13 and X30 and X51) xor (X13 and X31 and X50) xor (X13 and X31 and X51) xor (X13 and X31 and X53) xor (X13 and X33 and X50) xor (X20 and X30 and X51) xor (X20 and X31 and X50) xor (X20 and X31 and X53) xor (X20 and X33 and X51) xor (X20 and X33 and X53) xor (X21 and X30 and X51) xor (X21 and X30 and X53) xor (X21 and X31 and X53) xor (X21 and X33 and X50) xor (X21 and X33 and X51) xor (X21 and X33 and X53) xor (X23 and X30 and X51) xor (X23 and X31 and X50) xor (X23 and X31 and X51) xor (X23 and X31 and X53) xor (X23 and X33 and X50) xor (X43 and X53) xor (X43 and X50) xor (X43 and X51) xor (X41 and X50) xor (X00 and X40 and X51) xor (X00 and X41 and X50) xor (X00 and X41 and X53) xor (X00 and X43 and X51) xor (X00 and X43 and X53) xor (X0_1 and X40 and X51) xor (X0_1 and X40 and X53) xor (X0_1 and X41 and X53) xor (X0_1 and X43 and X50) xor (X0_1 and X43 and X51) xor (X0_1 and X43 and X53) xor (X03 and X40 and X51) xor (X03 and X41 and X50) xor (X03 and X41 and X51) xor (X03 and X41 and X53) xor (X03 and X43 and X50) xor (X10 and X40 and X51) xor (X10 and X41 and X50) xor (X10 and X41 and X53) xor (X10 and X43 and X51) xor (X10 and X43 and X53) xor (X11 and X40 and X51) xor (X11 and X40 and X53) xor (X11 and X41 and X53) xor (X11 and X43 and X50) xor (X11 and X43 and X51) xor (X11 and X43 and X53) xor (X13 and X40 and X51) xor (X13 and X41 and X50) xor (X13 and X41 and X51) xor (X13 and X41 and X53) xor (X13 and X43 and X50) xor (X03 and X63) xor (X03 and X60) xor (X03 and X61) xor (X0_1 and X60) xor (X13 and X63) xor (X13 and X60) xor (X13 and X61) xor (X11 and X60) xor (X00 and X20 and X61) xor (X00 and X21 and X60) xor (X00 and X21 and X63) xor (X00 and X23 and X61) xor (X00 and X23 and X63) xor (X0_1 and X20 and X61) xor (X0_1 and X20 and X63) xor (X0_1 and X21 and X63) xor (X0_1 and X23 and X60) xor (X0_1 and X23 and X61) xor (X0_1 and X23 and X63) xor (X03 and X20 and X61) xor (X03 and X21 and X60) xor (X03 and X21 and X61) xor (X03 and X21 and X63) xor (X03 and X23 and X60) xor (X33 and X63) xor (X33 and X60) xor (X33 and X61) xor (X31 and X60) xor (X20 and X30 and X61) xor (X20 and X31 and X60) xor (X20 and X31 and X63) xor (X20 and X33 and X61) xor (X20 and X33 and X63) xor (X21 and X30 and X61) xor (X21 and X30 and X63) xor (X21 and X31 and X63) xor (X21 and X33 and X60) xor (X21 and X33 and X61) xor (X21 and X33 and X63) xor (X23 and X30 and X61) xor (X23 and X31 and X60) xor (X23 and X31 and X61) xor (X23 and X31 and X63) xor (X23 and X33 and X60) xor (X00 and X40 and X61) xor (X00 and X41 and X60) xor (X00 and X41 and X63) xor (X00 and X43 and X61) xor (X00 and X43 and X63) xor (X0_1 and X40 and X61) xor (X0_1 and X40 and X63) xor (X0_1 and X41 and X63) xor (X0_1 and X43 and X60) xor (X0_1 and X43 and X61) xor (X0_1 and X43 and X63) xor (X03 and X40 and X61) xor (X03 and X41 and X60) xor (X03 and X41 and X61) xor (X03 and X41 and X63) xor (X03 and X43 and X60) xor (X10 and X40 and X61) xor (X10 and X41 and X60) xor (X10 and X41 and X63) xor (X10 and X43 and X61) xor (X10 and X43 and X63) xor (X11 and X40 and X61) xor (X11 and X40 and X63) xor (X11 and X41 and X63) xor (X11 and X43 and X60) xor (X11 and X43 and X61) xor (X11 and X43 and X63) xor (X13 and X40 and X61) xor (X13 and X41 and X60) xor (X13 and X41 and X61) xor (X13 and X41 and X63) xor (X13 and X43 and X60) xor (X53 and X63) xor (X53 and X60) xor (X53 and X61) xor (X51 and X60) xor (X00 and X50 and X61) xor (X00 and X51 and X60) xor (X00 and X51 and X63) xor (X00 and X53 and X61) xor (X00 and X53 and X63) xor (X0_1 and X50 and X61) xor (X0_1 and X50 and X63) xor (X0_1 and X51 and X63) xor (X0_1 and X53 and X60) xor (X0_1 and X53 and X61) xor (X0_1 and X53 and X63) xor (X03 and X50 and X61) xor (X03 and X51 and X60) xor (X03 and X51 and X61) xor (X03 and X51 and X63) xor (X03 and X53 and X60) xor (X40 and X50 and X61) xor (X40 and X51 and X60) xor (X40 and X51 and X63) xor (X40 and X53 and X61) xor (X40 and X53 and X63) xor (X41 and X50 and X61) xor (X41 and X50 and X63) xor (X41 and X51 and X63) xor (X41 and X53 and X60) xor (X41 and X53 and X61) xor (X41 and X53 and X63) xor (X43 and X50 and X61) xor (X43 and X51 and X60) xor (X43 and X51 and X61) xor (X43 and X51 and X63) xor (X43 and X53 and X60) xor (X73) xor (X03 and X73) xor (X03 and X70) xor (X03 and X71) xor (X0_1 and X70) xor (X13 and X73) xor (X13 and X70) xor (X13 and X71) xor (X11 and X70) xor (X00 and X10 and X71) xor (X00 and X11 and X70) xor (X00 and X11 and X73) xor (X00 and X13 and X71) xor (X00 and X13 and X73) xor (X0_1 and X10 and X71) xor (X0_1 and X10 and X73) xor (X0_1 and X11 and X73) xor (X0_1 and X13 and X70) xor (X0_1 and X13 and X71) xor (X0_1 and X13 and X73) xor (X03 and X10 and X71) xor (X03 and X11 and X70) xor (X03 and X11 and X71) xor (X03 and X11 and X73) xor (X03 and X13 and X70) xor (X23 and X73) xor (X23 and X70) xor (X23 and X71) xor (X21 and X70) xor (X43 and X73) xor (X43 and X70) xor (X43 and X71) xor (X41 and X70) xor (X00 and X40 and X71) xor (X00 and X41 and X70) xor (X00 and X41 and X73) xor (X00 and X43 and X71) xor (X00 and X43 and X73) xor (X0_1 and X40 and X71) xor (X0_1 and X40 and X73) xor (X0_1 and X41 and X73) xor (X0_1 and X43 and X70) xor (X0_1 and X43 and X71) xor (X0_1 and X43 and X73) xor (X03 and X40 and X71) xor (X03 and X41 and X70) xor (X03 and X41 and X71) xor (X03 and X41 and X73) xor (X03 and X43 and X70) xor (X53 and X73) xor (X53 and X70) xor (X53 and X71) xor (X51 and X70) xor (X00 and X50 and X71) xor (X00 and X51 and X70) xor (X00 and X51 and X73) xor (X00 and X53 and X71) xor (X00 and X53 and X73) xor (X0_1 and X50 and X71) xor (X0_1 and X50 and X73) xor (X0_1 and X51 and X73) xor (X0_1 and X53 and X70) xor (X0_1 and X53 and X71) xor (X0_1 and X53 and X73) xor (X03 and X50 and X71) xor (X03 and X51 and X70) xor (X03 and X51 and X71) xor (X03 and X51 and X73) xor (X03 and X53 and X70) xor (X20 and X50 and X71) xor (X20 and X51 and X70) xor (X20 and X51 and X73) xor (X20 and X53 and X71) xor (X20 and X53 and X73) xor (X21 and X50 and X71) xor (X21 and X50 and X73) xor (X21 and X51 and X73) xor (X21 and X53 and X70) xor (X21 and X53 and X71) xor (X21 and X53 and X73) xor (X23 and X50 and X71) xor (X23 and X51 and X70) xor (X23 and X51 and X71) xor (X23 and X51 and X73) xor (X23 and X53 and X70) xor (X40 and X50 and X71) xor (X40 and X51 and X70) xor (X40 and X51 and X73) xor (X40 and X53 and X71) xor (X40 and X53 and X73) xor (X41 and X50 and X71) xor (X41 and X50 and X73) xor (X41 and X51 and X73) xor (X41 and X53 and X70) xor (X41 and X53 and X71) xor (X41 and X53 and X73) xor (X43 and X50 and X71) xor (X43 and X51 and X70) xor (X43 and X51 and X71) xor (X43 and X51 and X73) xor (X43 and X53 and X70) xor (X20 and X60 and X71) xor (X20 and X61 and X70) xor (X20 and X61 and X73) xor (X20 and X63 and X71) xor (X20 and X63 and X73) xor (X21 and X60 and X71) xor (X21 and X60 and X73) xor (X21 and X61 and X73) xor (X21 and X63 and X70) xor (X21 and X63 and X71) xor (X21 and X63 and X73) xor (X23 and X60 and X71) xor (X23 and X61 and X70) xor (X23 and X61 and X71) xor (X23 and X61 and X73) xor (X23 and X63 and X70) xor (X30 and X60 and X71) xor (X30 and X61 and X70) xor (X30 and X61 and X73) xor (X30 and X63 and X71) xor (X30 and X63 and X73) xor (X31 and X60 and X71) xor (X31 and X60 and X73) xor (X31 and X61 and X73) xor (X31 and X63 and X70) xor (X31 and X63 and X71) xor (X31 and X63 and X73) xor (X33 and X60 and X71) xor (X33 and X61 and X70) xor (X33 and X61 and X71) xor (X33 and X61 and X73) xor (X33 and X63 and X70) xor (X40 and X60 and X71) xor (X40 and X61 and X70) xor (X40 and X61 and X73) xor (X40 and X63 and X71) xor (X40 and X63 and X73) xor (X41 and X60 and X71) xor (X41 and X60 and X73) xor (X41 and X61 and X73) xor (X41 and X63 and X70) xor (X41 and X63 and X71) xor (X41 and X63 and X73) xor (X43 and X60 and X71) xor (X43 and X61 and X70) xor (X43 and X61 and X71) xor (X43 and X61 and X73) xor (X43 and X63 and X70));
    F50  <= ((X00 and X10) xor (X00 and X11) xor (X02 and X10) xor (X00 and X12) xor (X20) xor (X00 and X20) xor (X00 and X21) xor (X02 and X20) xor (X00 and X22) xor (X00 and X30) xor (X00 and X31) xor (X02 and X30) xor (X00 and X32) xor (X00 and X10 and X30) xor (X00 and X10 and X32) xor (X00 and X11 and X31) xor (X00 and X11 and X32) xor (X00 and X12 and X31) xor (X0_1 and X10 and X30) xor (X0_1 and X10 and X32) xor (X0_1 and X11 and X30) xor (X0_1 and X12 and X30) xor (X0_1 and X12 and X31) xor (X02 and X10 and X30) xor (X02 and X10 and X31) xor (X02 and X11 and X30) xor (X02 and X11 and X31) xor (X02 and X12 and X30) xor (X02 and X12 and X32) xor (X00 and X40) xor (X00 and X41) xor (X02 and X40) xor (X00 and X42) xor (X20 and X40) xor (X20 and X41) xor (X22 and X40) xor (X20 and X42) xor (X00 and X20 and X40) xor (X00 and X20 and X42) xor (X00 and X21 and X41) xor (X00 and X21 and X42) xor (X00 and X22 and X41) xor (X0_1 and X20 and X40) xor (X0_1 and X20 and X42) xor (X0_1 and X21 and X40) xor (X0_1 and X22 and X40) xor (X0_1 and X22 and X41) xor (X02 and X20 and X40) xor (X02 and X20 and X41) xor (X02 and X21 and X40) xor (X02 and X21 and X41) xor (X02 and X22 and X40) xor (X02 and X22 and X42) xor (X10 and X20 and X40) xor (X10 and X20 and X42) xor (X10 and X21 and X41) xor (X10 and X21 and X42) xor (X10 and X22 and X41) xor (X11 and X20 and X40) xor (X11 and X20 and X42) xor (X11 and X21 and X40) xor (X11 and X22 and X40) xor (X11 and X22 and X41) xor (X12 and X20 and X40) xor (X12 and X20 and X41) xor (X12 and X21 and X40) xor (X12 and X21 and X41) xor (X12 and X22 and X40) xor (X12 and X22 and X42) xor (X30 and X40) xor (X30 and X41) xor (X32 and X40) xor (X30 and X42) xor (X50) xor (X00 and X50) xor (X00 and X51) xor (X02 and X50) xor (X00 and X52) xor (X00 and X10 and X50) xor (X00 and X10 and X52) xor (X00 and X11 and X51) xor (X00 and X11 and X52) xor (X00 and X12 and X51) xor (X0_1 and X10 and X50) xor (X0_1 and X10 and X52) xor (X0_1 and X11 and X50) xor (X0_1 and X12 and X50) xor (X0_1 and X12 and X51) xor (X02 and X10 and X50) xor (X02 and X10 and X51) xor (X02 and X11 and X50) xor (X02 and X11 and X51) xor (X02 and X12 and X50) xor (X02 and X12 and X52) xor (X20 and X50) xor (X20 and X51) xor (X22 and X50) xor (X20 and X52) xor (X30 and X50) xor (X30 and X51) xor (X32 and X50) xor (X30 and X52) xor (X10 and X30 and X50) xor (X10 and X30 and X52) xor (X10 and X31 and X51) xor (X10 and X31 and X52) xor (X10 and X32 and X51) xor (X11 and X30 and X50) xor (X11 and X30 and X52) xor (X11 and X31 and X50) xor (X11 and X32 and X50) xor (X11 and X32 and X51) xor (X12 and X30 and X50) xor (X12 and X30 and X51) xor (X12 and X31 and X50) xor (X12 and X31 and X51) xor (X12 and X32 and X50) xor (X12 and X32 and X52) xor (X40 and X50) xor (X40 and X51) xor (X42 and X50) xor (X40 and X52) xor (X10 and X60) xor (X10 and X61) xor (X12 and X60) xor (X10 and X62) xor (X00 and X20 and X60) xor (X00 and X20 and X62) xor (X00 and X21 and X61) xor (X00 and X21 and X62) xor (X00 and X22 and X61) xor (X0_1 and X20 and X60) xor (X0_1 and X20 and X62) xor (X0_1 and X21 and X60) xor (X0_1 and X22 and X60) xor (X0_1 and X22 and X61) xor (X02 and X20 and X60) xor (X02 and X20 and X61) xor (X02 and X21 and X60) xor (X02 and X21 and X61) xor (X02 and X22 and X60) xor (X02 and X22 and X62) xor (X30 and X60) xor (X30 and X61) xor (X32 and X60) xor (X30 and X62) xor (X10 and X30 and X60) xor (X10 and X30 and X62) xor (X10 and X31 and X61) xor (X10 and X31 and X62) xor (X10 and X32 and X61) xor (X11 and X30 and X60) xor (X11 and X30 and X62) xor (X11 and X31 and X60) xor (X11 and X32 and X60) xor (X11 and X32 and X61) xor (X12 and X30 and X60) xor (X12 and X30 and X61) xor (X12 and X31 and X60) xor (X12 and X31 and X61) xor (X12 and X32 and X60) xor (X12 and X32 and X62) xor (X40 and X60) xor (X40 and X61) xor (X42 and X60) xor (X40 and X62) xor (X00 and X40 and X60) xor (X00 and X40 and X62) xor (X00 and X41 and X61) xor (X00 and X41 and X62) xor (X00 and X42 and X61) xor (X0_1 and X40 and X60) xor (X0_1 and X40 and X62) xor (X0_1 and X41 and X60) xor (X0_1 and X42 and X60) xor (X0_1 and X42 and X61) xor (X02 and X40 and X60) xor (X02 and X40 and X61) xor (X02 and X41 and X60) xor (X02 and X41 and X61) xor (X02 and X42 and X60) xor (X02 and X42 and X62) xor (X10 and X40 and X60) xor (X10 and X40 and X62) xor (X10 and X41 and X61) xor (X10 and X41 and X62) xor (X10 and X42 and X61) xor (X11 and X40 and X60) xor (X11 and X40 and X62) xor (X11 and X41 and X60) xor (X11 and X42 and X60) xor (X11 and X42 and X61) xor (X12 and X40 and X60) xor (X12 and X40 and X61) xor (X12 and X41 and X60) xor (X12 and X41 and X61) xor (X12 and X42 and X60) xor (X12 and X42 and X62) xor (X20 and X40 and X60) xor (X20 and X40 and X62) xor (X20 and X41 and X61) xor (X20 and X41 and X62) xor (X20 and X42 and X61) xor (X21 and X40 and X60) xor (X21 and X40 and X62) xor (X21 and X41 and X60) xor (X21 and X42 and X60) xor (X21 and X42 and X61) xor (X22 and X40 and X60) xor (X22 and X40 and X61) xor (X22 and X41 and X60) xor (X22 and X41 and X61) xor (X22 and X42 and X60) xor (X22 and X42 and X62) xor (X50 and X60) xor (X50 and X61) xor (X52 and X60) xor (X50 and X62) xor (X10 and X50 and X60) xor (X10 and X50 and X62) xor (X10 and X51 and X61) xor (X10 and X51 and X62) xor (X10 and X52 and X61) xor (X11 and X50 and X60) xor (X11 and X50 and X62) xor (X11 and X51 and X60) xor (X11 and X52 and X60) xor (X11 and X52 and X61) xor (X12 and X50 and X60) xor (X12 and X50 and X61) xor (X12 and X51 and X60) xor (X12 and X51 and X61) xor (X12 and X52 and X60) xor (X12 and X52 and X62) xor (X20 and X50 and X60) xor (X20 and X50 and X62) xor (X20 and X51 and X61) xor (X20 and X51 and X62) xor (X20 and X52 and X61) xor (X21 and X50 and X60) xor (X21 and X50 and X62) xor (X21 and X51 and X60) xor (X21 and X52 and X60) xor (X21 and X52 and X61) xor (X22 and X50 and X60) xor (X22 and X50 and X61) xor (X22 and X51 and X60) xor (X22 and X51 and X61) xor (X22 and X52 and X60) xor (X22 and X52 and X62) xor (X40 and X50 and X60) xor (X40 and X50 and X62) xor (X40 and X51 and X61) xor (X40 and X51 and X62) xor (X40 and X52 and X61) xor (X41 and X50 and X60) xor (X41 and X50 and X62) xor (X41 and X51 and X60) xor (X41 and X52 and X60) xor (X41 and X52 and X61) xor (X42 and X50 and X60) xor (X42 and X50 and X61) xor (X42 and X51 and X60) xor (X42 and X51 and X61) xor (X42 and X52 and X60) xor (X42 and X52 and X62) xor (X10 and X70) xor (X10 and X71) xor (X12 and X70) xor (X10 and X72) xor (X20 and X70) xor (X20 and X71) xor (X22 and X70) xor (X20 and X72) xor (X30 and X70) xor (X30 and X71) xor (X32 and X70) xor (X30 and X72) xor (X00 and X30 and X70) xor (X00 and X30 and X72) xor (X00 and X31 and X71) xor (X00 and X31 and X72) xor (X00 and X32 and X71) xor (X0_1 and X30 and X70) xor (X0_1 and X30 and X72) xor (X0_1 and X31 and X70) xor (X0_1 and X32 and X70) xor (X0_1 and X32 and X71) xor (X02 and X30 and X70) xor (X02 and X30 and X71) xor (X02 and X31 and X70) xor (X02 and X31 and X71) xor (X02 and X32 and X70) xor (X02 and X32 and X72) xor (X10 and X30 and X70) xor (X10 and X30 and X72) xor (X10 and X31 and X71) xor (X10 and X31 and X72) xor (X10 and X32 and X71) xor (X11 and X30 and X70) xor (X11 and X30 and X72) xor (X11 and X31 and X70) xor (X11 and X32 and X70) xor (X11 and X32 and X71) xor (X12 and X30 and X70) xor (X12 and X30 and X71) xor (X12 and X31 and X70) xor (X12 and X31 and X71) xor (X12 and X32 and X70) xor (X12 and X32 and X72) xor (X00 and X40 and X70) xor (X00 and X40 and X72) xor (X00 and X41 and X71) xor (X00 and X41 and X72) xor (X00 and X42 and X71) xor (X0_1 and X40 and X70) xor (X0_1 and X40 and X72) xor (X0_1 and X41 and X70) xor (X0_1 and X42 and X70) xor (X0_1 and X42 and X71) xor (X02 and X40 and X70) xor (X02 and X40 and X71) xor (X02 and X41 and X70) xor (X02 and X41 and X71) xor (X02 and X42 and X70) xor (X02 and X42 and X72) xor (X00 and X50 and X70) xor (X00 and X50 and X72) xor (X00 and X51 and X71) xor (X00 and X51 and X72) xor (X00 and X52 and X71) xor (X0_1 and X50 and X70) xor (X0_1 and X50 and X72) xor (X0_1 and X51 and X70) xor (X0_1 and X52 and X70) xor (X0_1 and X52 and X71) xor (X02 and X50 and X70) xor (X02 and X50 and X71) xor (X02 and X51 and X70) xor (X02 and X51 and X71) xor (X02 and X52 and X70) xor (X02 and X52 and X72) xor (X10 and X50 and X70) xor (X10 and X50 and X72) xor (X10 and X51 and X71) xor (X10 and X51 and X72) xor (X10 and X52 and X71) xor (X11 and X50 and X70) xor (X11 and X50 and X72) xor (X11 and X51 and X70) xor (X11 and X52 and X70) xor (X11 and X52 and X71) xor (X12 and X50 and X70) xor (X12 and X50 and X71) xor (X12 and X51 and X70) xor (X12 and X51 and X71) xor (X12 and X52 and X70) xor (X12 and X52 and X72) xor (X20 and X50 and X70) xor (X20 and X50 and X72) xor (X20 and X51 and X71) xor (X20 and X51 and X72) xor (X20 and X52 and X71) xor (X21 and X50 and X70) xor (X21 and X50 and X72) xor (X21 and X51 and X70) xor (X21 and X52 and X70) xor (X21 and X52 and X71) xor (X22 and X50 and X70) xor (X22 and X50 and X71) xor (X22 and X51 and X70) xor (X22 and X51 and X71) xor (X22 and X52 and X70) xor (X22 and X52 and X72) xor (X30 and X50 and X70) xor (X30 and X50 and X72) xor (X30 and X51 and X71) xor (X30 and X51 and X72) xor (X30 and X52 and X71) xor (X31 and X50 and X70) xor (X31 and X50 and X72) xor (X31 and X51 and X70) xor (X31 and X52 and X70) xor (X31 and X52 and X71) xor (X32 and X50 and X70) xor (X32 and X50 and X71) xor (X32 and X51 and X70) xor (X32 and X51 and X71) xor (X32 and X52 and X70) xor (X32 and X52 and X72) xor (X10 and X60 and X70) xor (X10 and X60 and X72) xor (X10 and X61 and X71) xor (X10 and X61 and X72) xor (X10 and X62 and X71) xor (X11 and X60 and X70) xor (X11 and X60 and X72) xor (X11 and X61 and X70) xor (X11 and X62 and X70) xor (X11 and X62 and X71) xor (X12 and X60 and X70) xor (X12 and X60 and X71) xor (X12 and X61 and X70) xor (X12 and X61 and X71) xor (X12 and X62 and X70) xor (X12 and X62 and X72) xor (X20 and X60 and X70) xor (X20 and X60 and X72) xor (X20 and X61 and X71) xor (X20 and X61 and X72) xor (X20 and X62 and X71) xor (X21 and X60 and X70) xor (X21 and X60 and X72) xor (X21 and X61 and X70) xor (X21 and X62 and X70) xor (X21 and X62 and X71) xor (X22 and X60 and X70) xor (X22 and X60 and X71) xor (X22 and X61 and X70) xor (X22 and X61 and X71) xor (X22 and X62 and X70) xor (X22 and X62 and X72) xor (X30 and X60 and X70) xor (X30 and X60 and X72) xor (X30 and X61 and X71) xor (X30 and X61 and X72) xor (X30 and X62 and X71) xor (X31 and X60 and X70) xor (X31 and X60 and X72) xor (X31 and X61 and X70) xor (X31 and X62 and X70) xor (X31 and X62 and X71) xor (X32 and X60 and X70) xor (X32 and X60 and X71) xor (X32 and X61 and X70) xor (X32 and X61 and X71) xor (X32 and X62 and X70) xor (X32 and X62 and X72) xor (X40 and X60 and X70) xor (X40 and X60 and X72) xor (X40 and X61 and X71) xor (X40 and X61 and X72) xor (X40 and X62 and X71) xor (X41 and X60 and X70) xor (X41 and X60 and X72) xor (X41 and X61 and X70) xor (X41 and X62 and X70) xor (X41 and X62 and X71) xor (X42 and X60 and X70) xor (X42 and X60 and X71) xor (X42 and X61 and X70) xor (X42 and X61 and X71) xor (X42 and X62 and X70) xor (X42 and X62 and X72) xor (X50 and X60 and X70) xor (X50 and X60 and X72) xor (X50 and X61 and X71) xor (X50 and X61 and X72) xor (X50 and X62 and X71) xor (X51 and X60 and X70) xor (X51 and X60 and X72) xor (X51 and X61 and X70) xor (X51 and X62 and X70) xor (X51 and X62 and X71) xor (X52 and X60 and X70) xor (X52 and X60 and X71) xor (X52 and X61 and X70) xor (X52 and X61 and X71) xor (X52 and X62 and X70) xor (X52 and X62 and X72));
    F51  <= ((X0_1 and X11) xor (X0_1 and X12) xor (X02 and X11) xor (X0_1 and X13) xor (X21) xor (X0_1 and X21) xor (X0_1 and X22) xor (X02 and X21) xor (X0_1 and X23) xor (X0_1 and X31) xor (X0_1 and X32) xor (X02 and X31) xor (X0_1 and X33) xor (X0_1 and X11 and X31) xor (X0_1 and X11 and X32) xor (X0_1 and X12 and X32) xor (X0_1 and X12 and X33) xor (X0_1 and X13 and X32) xor (X02 and X11 and X32) xor (X02 and X11 and X33) xor (X02 and X12 and X31) xor (X02 and X12 and X33) xor (X02 and X13 and X31) xor (X02 and X13 and X32) xor (X03 and X11 and X32) xor (X03 and X12 and X31) xor (X03 and X12 and X33) xor (X03 and X13 and X31) xor (X03 and X13 and X33) xor (X0_1 and X41) xor (X0_1 and X42) xor (X02 and X41) xor (X0_1 and X43) xor (X21 and X41) xor (X21 and X42) xor (X22 and X41) xor (X21 and X43) xor (X0_1 and X21 and X41) xor (X0_1 and X21 and X42) xor (X0_1 and X22 and X42) xor (X0_1 and X22 and X43) xor (X0_1 and X23 and X42) xor (X02 and X21 and X42) xor (X02 and X21 and X43) xor (X02 and X22 and X41) xor (X02 and X22 and X43) xor (X02 and X23 and X41) xor (X02 and X23 and X42) xor (X03 and X21 and X42) xor (X03 and X22 and X41) xor (X03 and X22 and X43) xor (X03 and X23 and X41) xor (X03 and X23 and X43) xor (X11 and X21 and X41) xor (X11 and X21 and X42) xor (X11 and X22 and X42) xor (X11 and X22 and X43) xor (X11 and X23 and X42) xor (X12 and X21 and X42) xor (X12 and X21 and X43) xor (X12 and X22 and X41) xor (X12 and X22 and X43) xor (X12 and X23 and X41) xor (X12 and X23 and X42) xor (X13 and X21 and X42) xor (X13 and X22 and X41) xor (X13 and X22 and X43) xor (X13 and X23 and X41) xor (X13 and X23 and X43) xor (X31 and X41) xor (X31 and X42) xor (X32 and X41) xor (X31 and X43) xor (X51) xor (X0_1 and X51) xor (X0_1 and X52) xor (X02 and X51) xor (X0_1 and X53) xor (X0_1 and X11 and X51) xor (X0_1 and X11 and X52) xor (X0_1 and X12 and X52) xor (X0_1 and X12 and X53) xor (X0_1 and X13 and X52) xor (X02 and X11 and X52) xor (X02 and X11 and X53) xor (X02 and X12 and X51) xor (X02 and X12 and X53) xor (X02 and X13 and X51) xor (X02 and X13 and X52) xor (X03 and X11 and X52) xor (X03 and X12 and X51) xor (X03 and X12 and X53) xor (X03 and X13 and X51) xor (X03 and X13 and X53) xor (X21 and X51) xor (X21 and X52) xor (X22 and X51) xor (X21 and X53) xor (X31 and X51) xor (X31 and X52) xor (X32 and X51) xor (X31 and X53) xor (X11 and X31 and X51) xor (X11 and X31 and X52) xor (X11 and X32 and X52) xor (X11 and X32 and X53) xor (X11 and X33 and X52) xor (X12 and X31 and X52) xor (X12 and X31 and X53) xor (X12 and X32 and X51) xor (X12 and X32 and X53) xor (X12 and X33 and X51) xor (X12 and X33 and X52) xor (X13 and X31 and X52) xor (X13 and X32 and X51) xor (X13 and X32 and X53) xor (X13 and X33 and X51) xor (X13 and X33 and X53) xor (X41 and X51) xor (X41 and X52) xor (X42 and X51) xor (X41 and X53) xor (X11 and X61) xor (X11 and X62) xor (X12 and X61) xor (X11 and X63) xor (X0_1 and X21 and X61) xor (X0_1 and X21 and X62) xor (X0_1 and X22 and X62) xor (X0_1 and X22 and X63) xor (X0_1 and X23 and X62) xor (X02 and X21 and X62) xor (X02 and X21 and X63) xor (X02 and X22 and X61) xor (X02 and X22 and X63) xor (X02 and X23 and X61) xor (X02 and X23 and X62) xor (X03 and X21 and X62) xor (X03 and X22 and X61) xor (X03 and X22 and X63) xor (X03 and X23 and X61) xor (X03 and X23 and X63) xor (X31 and X61) xor (X31 and X62) xor (X32 and X61) xor (X31 and X63) xor (X11 and X31 and X61) xor (X11 and X31 and X62) xor (X11 and X32 and X62) xor (X11 and X32 and X63) xor (X11 and X33 and X62) xor (X12 and X31 and X62) xor (X12 and X31 and X63) xor (X12 and X32 and X61) xor (X12 and X32 and X63) xor (X12 and X33 and X61) xor (X12 and X33 and X62) xor (X13 and X31 and X62) xor (X13 and X32 and X61) xor (X13 and X32 and X63) xor (X13 and X33 and X61) xor (X13 and X33 and X63) xor (X41 and X61) xor (X41 and X62) xor (X42 and X61) xor (X41 and X63) xor (X0_1 and X41 and X61) xor (X0_1 and X41 and X62) xor (X0_1 and X42 and X62) xor (X0_1 and X42 and X63) xor (X0_1 and X43 and X62) xor (X02 and X41 and X62) xor (X02 and X41 and X63) xor (X02 and X42 and X61) xor (X02 and X42 and X63) xor (X02 and X43 and X61) xor (X02 and X43 and X62) xor (X03 and X41 and X62) xor (X03 and X42 and X61) xor (X03 and X42 and X63) xor (X03 and X43 and X61) xor (X03 and X43 and X63) xor (X11 and X41 and X61) xor (X11 and X41 and X62) xor (X11 and X42 and X62) xor (X11 and X42 and X63) xor (X11 and X43 and X62) xor (X12 and X41 and X62) xor (X12 and X41 and X63) xor (X12 and X42 and X61) xor (X12 and X42 and X63) xor (X12 and X43 and X61) xor (X12 and X43 and X62) xor (X13 and X41 and X62) xor (X13 and X42 and X61) xor (X13 and X42 and X63) xor (X13 and X43 and X61) xor (X13 and X43 and X63) xor (X21 and X41 and X61) xor (X21 and X41 and X62) xor (X21 and X42 and X62) xor (X21 and X42 and X63) xor (X21 and X43 and X62) xor (X22 and X41 and X62) xor (X22 and X41 and X63) xor (X22 and X42 and X61) xor (X22 and X42 and X63) xor (X22 and X43 and X61) xor (X22 and X43 and X62) xor (X23 and X41 and X62) xor (X23 and X42 and X61) xor (X23 and X42 and X63) xor (X23 and X43 and X61) xor (X23 and X43 and X63) xor (X51 and X61) xor (X51 and X62) xor (X52 and X61) xor (X51 and X63) xor (X11 and X51 and X61) xor (X11 and X51 and X62) xor (X11 and X52 and X62) xor (X11 and X52 and X63) xor (X11 and X53 and X62) xor (X12 and X51 and X62) xor (X12 and X51 and X63) xor (X12 and X52 and X61) xor (X12 and X52 and X63) xor (X12 and X53 and X61) xor (X12 and X53 and X62) xor (X13 and X51 and X62) xor (X13 and X52 and X61) xor (X13 and X52 and X63) xor (X13 and X53 and X61) xor (X13 and X53 and X63) xor (X21 and X51 and X61) xor (X21 and X51 and X62) xor (X21 and X52 and X62) xor (X21 and X52 and X63) xor (X21 and X53 and X62) xor (X22 and X51 and X62) xor (X22 and X51 and X63) xor (X22 and X52 and X61) xor (X22 and X52 and X63) xor (X22 and X53 and X61) xor (X22 and X53 and X62) xor (X23 and X51 and X62) xor (X23 and X52 and X61) xor (X23 and X52 and X63) xor (X23 and X53 and X61) xor (X23 and X53 and X63) xor (X41 and X51 and X61) xor (X41 and X51 and X62) xor (X41 and X52 and X62) xor (X41 and X52 and X63) xor (X41 and X53 and X62) xor (X42 and X51 and X62) xor (X42 and X51 and X63) xor (X42 and X52 and X61) xor (X42 and X52 and X63) xor (X42 and X53 and X61) xor (X42 and X53 and X62) xor (X43 and X51 and X62) xor (X43 and X52 and X61) xor (X43 and X52 and X63) xor (X43 and X53 and X61) xor (X43 and X53 and X63) xor (X11 and X71) xor (X11 and X72) xor (X12 and X71) xor (X11 and X73) xor (X21 and X71) xor (X21 and X72) xor (X22 and X71) xor (X21 and X73) xor (X31 and X71) xor (X31 and X72) xor (X32 and X71) xor (X31 and X73) xor (X0_1 and X31 and X71) xor (X0_1 and X31 and X72) xor (X0_1 and X32 and X72) xor (X0_1 and X32 and X73) xor (X0_1 and X33 and X72) xor (X02 and X31 and X72) xor (X02 and X31 and X73) xor (X02 and X32 and X71) xor (X02 and X32 and X73) xor (X02 and X33 and X71) xor (X02 and X33 and X72) xor (X03 and X31 and X72) xor (X03 and X32 and X71) xor (X03 and X32 and X73) xor (X03 and X33 and X71) xor (X03 and X33 and X73) xor (X11 and X31 and X71) xor (X11 and X31 and X72) xor (X11 and X32 and X72) xor (X11 and X32 and X73) xor (X11 and X33 and X72) xor (X12 and X31 and X72) xor (X12 and X31 and X73) xor (X12 and X32 and X71) xor (X12 and X32 and X73) xor (X12 and X33 and X71) xor (X12 and X33 and X72) xor (X13 and X31 and X72) xor (X13 and X32 and X71) xor (X13 and X32 and X73) xor (X13 and X33 and X71) xor (X13 and X33 and X73) xor (X0_1 and X41 and X71) xor (X0_1 and X41 and X72) xor (X0_1 and X42 and X72) xor (X0_1 and X42 and X73) xor (X0_1 and X43 and X72) xor (X02 and X41 and X72) xor (X02 and X41 and X73) xor (X02 and X42 and X71) xor (X02 and X42 and X73) xor (X02 and X43 and X71) xor (X02 and X43 and X72) xor (X03 and X41 and X72) xor (X03 and X42 and X71) xor (X03 and X42 and X73) xor (X03 and X43 and X71) xor (X03 and X43 and X73) xor (X0_1 and X51 and X71) xor (X0_1 and X51 and X72) xor (X0_1 and X52 and X72) xor (X0_1 and X52 and X73) xor (X0_1 and X53 and X72) xor (X02 and X51 and X72) xor (X02 and X51 and X73) xor (X02 and X52 and X71) xor (X02 and X52 and X73) xor (X02 and X53 and X71) xor (X02 and X53 and X72) xor (X03 and X51 and X72) xor (X03 and X52 and X71) xor (X03 and X52 and X73) xor (X03 and X53 and X71) xor (X03 and X53 and X73) xor (X11 and X51 and X71) xor (X11 and X51 and X72) xor (X11 and X52 and X72) xor (X11 and X52 and X73) xor (X11 and X53 and X72) xor (X12 and X51 and X72) xor (X12 and X51 and X73) xor (X12 and X52 and X71) xor (X12 and X52 and X73) xor (X12 and X53 and X71) xor (X12 and X53 and X72) xor (X13 and X51 and X72) xor (X13 and X52 and X71) xor (X13 and X52 and X73) xor (X13 and X53 and X71) xor (X13 and X53 and X73) xor (X21 and X51 and X71) xor (X21 and X51 and X72) xor (X21 and X52 and X72) xor (X21 and X52 and X73) xor (X21 and X53 and X72) xor (X22 and X51 and X72) xor (X22 and X51 and X73) xor (X22 and X52 and X71) xor (X22 and X52 and X73) xor (X22 and X53 and X71) xor (X22 and X53 and X72) xor (X23 and X51 and X72) xor (X23 and X52 and X71) xor (X23 and X52 and X73) xor (X23 and X53 and X71) xor (X23 and X53 and X73) xor (X31 and X51 and X71) xor (X31 and X51 and X72) xor (X31 and X52 and X72) xor (X31 and X52 and X73) xor (X31 and X53 and X72) xor (X32 and X51 and X72) xor (X32 and X51 and X73) xor (X32 and X52 and X71) xor (X32 and X52 and X73) xor (X32 and X53 and X71) xor (X32 and X53 and X72) xor (X33 and X51 and X72) xor (X33 and X52 and X71) xor (X33 and X52 and X73) xor (X33 and X53 and X71) xor (X33 and X53 and X73) xor (X11 and X61 and X71) xor (X11 and X61 and X72) xor (X11 and X62 and X72) xor (X11 and X62 and X73) xor (X11 and X63 and X72) xor (X12 and X61 and X72) xor (X12 and X61 and X73) xor (X12 and X62 and X71) xor (X12 and X62 and X73) xor (X12 and X63 and X71) xor (X12 and X63 and X72) xor (X13 and X61 and X72) xor (X13 and X62 and X71) xor (X13 and X62 and X73) xor (X13 and X63 and X71) xor (X13 and X63 and X73) xor (X21 and X61 and X71) xor (X21 and X61 and X72) xor (X21 and X62 and X72) xor (X21 and X62 and X73) xor (X21 and X63 and X72) xor (X22 and X61 and X72) xor (X22 and X61 and X73) xor (X22 and X62 and X71) xor (X22 and X62 and X73) xor (X22 and X63 and X71) xor (X22 and X63 and X72) xor (X23 and X61 and X72) xor (X23 and X62 and X71) xor (X23 and X62 and X73) xor (X23 and X63 and X71) xor (X23 and X63 and X73) xor (X31 and X61 and X71) xor (X31 and X61 and X72) xor (X31 and X62 and X72) xor (X31 and X62 and X73) xor (X31 and X63 and X72) xor (X32 and X61 and X72) xor (X32 and X61 and X73) xor (X32 and X62 and X71) xor (X32 and X62 and X73) xor (X32 and X63 and X71) xor (X32 and X63 and X72) xor (X33 and X61 and X72) xor (X33 and X62 and X71) xor (X33 and X62 and X73) xor (X33 and X63 and X71) xor (X33 and X63 and X73) xor (X41 and X61 and X71) xor (X41 and X61 and X72) xor (X41 and X62 and X72) xor (X41 and X62 and X73) xor (X41 and X63 and X72) xor (X42 and X61 and X72) xor (X42 and X61 and X73) xor (X42 and X62 and X71) xor (X42 and X62 and X73) xor (X42 and X63 and X71) xor (X42 and X63 and X72) xor (X43 and X61 and X72) xor (X43 and X62 and X71) xor (X43 and X62 and X73) xor (X43 and X63 and X71) xor (X43 and X63 and X73) xor (X51 and X61 and X71) xor (X51 and X61 and X72) xor (X51 and X62 and X72) xor (X51 and X62 and X73) xor (X51 and X63 and X72) xor (X52 and X61 and X72) xor (X52 and X61 and X73) xor (X52 and X62 and X71) xor (X52 and X62 and X73) xor (X52 and X63 and X71) xor (X52 and X63 and X72) xor (X53 and X61 and X72) xor (X53 and X62 and X71) xor (X53 and X62 and X73) xor (X53 and X63 and X71) xor (X53 and X63 and X73));
    F52  <= ((X02 and X12) xor (X00 and X13) xor (X02 and X13) xor (X03 and X12) xor (X22) xor (X02 and X22) xor (X00 and X23) xor (X02 and X23) xor (X03 and X22) xor (X02 and X32) xor (X00 and X33) xor (X02 and X33) xor (X03 and X32) xor (X00 and X10 and X33) xor (X00 and X12 and X30) xor (X00 and X12 and X32) xor (X00 and X12 and X33) xor (X00 and X13 and X30) xor (X00 and X13 and X32) xor (X02 and X10 and X32) xor (X02 and X10 and X33) xor (X02 and X13 and X30) xor (X02 and X13 and X33) xor (X03 and X10 and X30) xor (X03 and X10 and X32) xor (X03 and X10 and X33) xor (X03 and X12 and X30) xor (X03 and X12 and X32) xor (X03 and X13 and X32) xor (X02 and X42) xor (X00 and X43) xor (X02 and X43) xor (X03 and X42) xor (X22 and X42) xor (X20 and X43) xor (X22 and X43) xor (X23 and X42) xor (X00 and X20 and X43) xor (X00 and X22 and X40) xor (X00 and X22 and X42) xor (X00 and X22 and X43) xor (X00 and X23 and X40) xor (X00 and X23 and X42) xor (X02 and X20 and X42) xor (X02 and X20 and X43) xor (X02 and X23 and X40) xor (X02 and X23 and X43) xor (X03 and X20 and X40) xor (X03 and X20 and X42) xor (X03 and X20 and X43) xor (X03 and X22 and X40) xor (X03 and X22 and X42) xor (X03 and X23 and X42) xor (X10 and X20 and X43) xor (X10 and X22 and X40) xor (X10 and X22 and X42) xor (X10 and X22 and X43) xor (X10 and X23 and X40) xor (X10 and X23 and X42) xor (X12 and X20 and X42) xor (X12 and X20 and X43) xor (X12 and X23 and X40) xor (X12 and X23 and X43) xor (X13 and X20 and X40) xor (X13 and X20 and X42) xor (X13 and X20 and X43) xor (X13 and X22 and X40) xor (X13 and X22 and X42) xor (X13 and X23 and X42) xor (X32 and X42) xor (X30 and X43) xor (X32 and X43) xor (X33 and X42) xor (X52) xor (X02 and X52) xor (X00 and X53) xor (X02 and X53) xor (X03 and X52) xor (X00 and X10 and X53) xor (X00 and X12 and X50) xor (X00 and X12 and X52) xor (X00 and X12 and X53) xor (X00 and X13 and X50) xor (X00 and X13 and X52) xor (X02 and X10 and X52) xor (X02 and X10 and X53) xor (X02 and X13 and X50) xor (X02 and X13 and X53) xor (X03 and X10 and X50) xor (X03 and X10 and X52) xor (X03 and X10 and X53) xor (X03 and X12 and X50) xor (X03 and X12 and X52) xor (X03 and X13 and X52) xor (X22 and X52) xor (X20 and X53) xor (X22 and X53) xor (X23 and X52) xor (X32 and X52) xor (X30 and X53) xor (X32 and X53) xor (X33 and X52) xor (X10 and X30 and X53) xor (X10 and X32 and X50) xor (X10 and X32 and X52) xor (X10 and X32 and X53) xor (X10 and X33 and X50) xor (X10 and X33 and X52) xor (X12 and X30 and X52) xor (X12 and X30 and X53) xor (X12 and X33 and X50) xor (X12 and X33 and X53) xor (X13 and X30 and X50) xor (X13 and X30 and X52) xor (X13 and X30 and X53) xor (X13 and X32 and X50) xor (X13 and X32 and X52) xor (X13 and X33 and X52) xor (X42 and X52) xor (X40 and X53) xor (X42 and X53) xor (X43 and X52) xor (X12 and X62) xor (X10 and X63) xor (X12 and X63) xor (X13 and X62) xor (X00 and X20 and X63) xor (X00 and X22 and X60) xor (X00 and X22 and X62) xor (X00 and X22 and X63) xor (X00 and X23 and X60) xor (X00 and X23 and X62) xor (X02 and X20 and X62) xor (X02 and X20 and X63) xor (X02 and X23 and X60) xor (X02 and X23 and X63) xor (X03 and X20 and X60) xor (X03 and X20 and X62) xor (X03 and X20 and X63) xor (X03 and X22 and X60) xor (X03 and X22 and X62) xor (X03 and X23 and X62) xor (X32 and X62) xor (X30 and X63) xor (X32 and X63) xor (X33 and X62) xor (X10 and X30 and X63) xor (X10 and X32 and X60) xor (X10 and X32 and X62) xor (X10 and X32 and X63) xor (X10 and X33 and X60) xor (X10 and X33 and X62) xor (X12 and X30 and X62) xor (X12 and X30 and X63) xor (X12 and X33 and X60) xor (X12 and X33 and X63) xor (X13 and X30 and X60) xor (X13 and X30 and X62) xor (X13 and X30 and X63) xor (X13 and X32 and X60) xor (X13 and X32 and X62) xor (X13 and X33 and X62) xor (X42 and X62) xor (X40 and X63) xor (X42 and X63) xor (X43 and X62) xor (X00 and X40 and X63) xor (X00 and X42 and X60) xor (X00 and X42 and X62) xor (X00 and X42 and X63) xor (X00 and X43 and X60) xor (X00 and X43 and X62) xor (X02 and X40 and X62) xor (X02 and X40 and X63) xor (X02 and X43 and X60) xor (X02 and X43 and X63) xor (X03 and X40 and X60) xor (X03 and X40 and X62) xor (X03 and X40 and X63) xor (X03 and X42 and X60) xor (X03 and X42 and X62) xor (X03 and X43 and X62) xor (X10 and X40 and X63) xor (X10 and X42 and X60) xor (X10 and X42 and X62) xor (X10 and X42 and X63) xor (X10 and X43 and X60) xor (X10 and X43 and X62) xor (X12 and X40 and X62) xor (X12 and X40 and X63) xor (X12 and X43 and X60) xor (X12 and X43 and X63) xor (X13 and X40 and X60) xor (X13 and X40 and X62) xor (X13 and X40 and X63) xor (X13 and X42 and X60) xor (X13 and X42 and X62) xor (X13 and X43 and X62) xor (X20 and X40 and X63) xor (X20 and X42 and X60) xor (X20 and X42 and X62) xor (X20 and X42 and X63) xor (X20 and X43 and X60) xor (X20 and X43 and X62) xor (X22 and X40 and X62) xor (X22 and X40 and X63) xor (X22 and X43 and X60) xor (X22 and X43 and X63) xor (X23 and X40 and X60) xor (X23 and X40 and X62) xor (X23 and X40 and X63) xor (X23 and X42 and X60) xor (X23 and X42 and X62) xor (X23 and X43 and X62) xor (X52 and X62) xor (X50 and X63) xor (X52 and X63) xor (X53 and X62) xor (X10 and X50 and X63) xor (X10 and X52 and X60) xor (X10 and X52 and X62) xor (X10 and X52 and X63) xor (X10 and X53 and X60) xor (X10 and X53 and X62) xor (X12 and X50 and X62) xor (X12 and X50 and X63) xor (X12 and X53 and X60) xor (X12 and X53 and X63) xor (X13 and X50 and X60) xor (X13 and X50 and X62) xor (X13 and X50 and X63) xor (X13 and X52 and X60) xor (X13 and X52 and X62) xor (X13 and X53 and X62) xor (X20 and X50 and X63) xor (X20 and X52 and X60) xor (X20 and X52 and X62) xor (X20 and X52 and X63) xor (X20 and X53 and X60) xor (X20 and X53 and X62) xor (X22 and X50 and X62) xor (X22 and X50 and X63) xor (X22 and X53 and X60) xor (X22 and X53 and X63) xor (X23 and X50 and X60) xor (X23 and X50 and X62) xor (X23 and X50 and X63) xor (X23 and X52 and X60) xor (X23 and X52 and X62) xor (X23 and X53 and X62) xor (X40 and X50 and X63) xor (X40 and X52 and X60) xor (X40 and X52 and X62) xor (X40 and X52 and X63) xor (X40 and X53 and X60) xor (X40 and X53 and X62) xor (X42 and X50 and X62) xor (X42 and X50 and X63) xor (X42 and X53 and X60) xor (X42 and X53 and X63) xor (X43 and X50 and X60) xor (X43 and X50 and X62) xor (X43 and X50 and X63) xor (X43 and X52 and X60) xor (X43 and X52 and X62) xor (X43 and X53 and X62) xor (X12 and X72) xor (X10 and X73) xor (X12 and X73) xor (X13 and X72) xor (X22 and X72) xor (X20 and X73) xor (X22 and X73) xor (X23 and X72) xor (X32 and X72) xor (X30 and X73) xor (X32 and X73) xor (X33 and X72) xor (X00 and X30 and X73) xor (X00 and X32 and X70) xor (X00 and X32 and X72) xor (X00 and X32 and X73) xor (X00 and X33 and X70) xor (X00 and X33 and X72) xor (X02 and X30 and X72) xor (X02 and X30 and X73) xor (X02 and X33 and X70) xor (X02 and X33 and X73) xor (X03 and X30 and X70) xor (X03 and X30 and X72) xor (X03 and X30 and X73) xor (X03 and X32 and X70) xor (X03 and X32 and X72) xor (X03 and X33 and X72) xor (X10 and X30 and X73) xor (X10 and X32 and X70) xor (X10 and X32 and X72) xor (X10 and X32 and X73) xor (X10 and X33 and X70) xor (X10 and X33 and X72) xor (X12 and X30 and X72) xor (X12 and X30 and X73) xor (X12 and X33 and X70) xor (X12 and X33 and X73) xor (X13 and X30 and X70) xor (X13 and X30 and X72) xor (X13 and X30 and X73) xor (X13 and X32 and X70) xor (X13 and X32 and X72) xor (X13 and X33 and X72) xor (X00 and X40 and X73) xor (X00 and X42 and X70) xor (X00 and X42 and X72) xor (X00 and X42 and X73) xor (X00 and X43 and X70) xor (X00 and X43 and X72) xor (X02 and X40 and X72) xor (X02 and X40 and X73) xor (X02 and X43 and X70) xor (X02 and X43 and X73) xor (X03 and X40 and X70) xor (X03 and X40 and X72) xor (X03 and X40 and X73) xor (X03 and X42 and X70) xor (X03 and X42 and X72) xor (X03 and X43 and X72) xor (X00 and X50 and X73) xor (X00 and X52 and X70) xor (X00 and X52 and X72) xor (X00 and X52 and X73) xor (X00 and X53 and X70) xor (X00 and X53 and X72) xor (X02 and X50 and X72) xor (X02 and X50 and X73) xor (X02 and X53 and X70) xor (X02 and X53 and X73) xor (X03 and X50 and X70) xor (X03 and X50 and X72) xor (X03 and X50 and X73) xor (X03 and X52 and X70) xor (X03 and X52 and X72) xor (X03 and X53 and X72) xor (X10 and X50 and X73) xor (X10 and X52 and X70) xor (X10 and X52 and X72) xor (X10 and X52 and X73) xor (X10 and X53 and X70) xor (X10 and X53 and X72) xor (X12 and X50 and X72) xor (X12 and X50 and X73) xor (X12 and X53 and X70) xor (X12 and X53 and X73) xor (X13 and X50 and X70) xor (X13 and X50 and X72) xor (X13 and X50 and X73) xor (X13 and X52 and X70) xor (X13 and X52 and X72) xor (X13 and X53 and X72) xor (X20 and X50 and X73) xor (X20 and X52 and X70) xor (X20 and X52 and X72) xor (X20 and X52 and X73) xor (X20 and X53 and X70) xor (X20 and X53 and X72) xor (X22 and X50 and X72) xor (X22 and X50 and X73) xor (X22 and X53 and X70) xor (X22 and X53 and X73) xor (X23 and X50 and X70) xor (X23 and X50 and X72) xor (X23 and X50 and X73) xor (X23 and X52 and X70) xor (X23 and X52 and X72) xor (X23 and X53 and X72) xor (X30 and X50 and X73) xor (X30 and X52 and X70) xor (X30 and X52 and X72) xor (X30 and X52 and X73) xor (X30 and X53 and X70) xor (X30 and X53 and X72) xor (X32 and X50 and X72) xor (X32 and X50 and X73) xor (X32 and X53 and X70) xor (X32 and X53 and X73) xor (X33 and X50 and X70) xor (X33 and X50 and X72) xor (X33 and X50 and X73) xor (X33 and X52 and X70) xor (X33 and X52 and X72) xor (X33 and X53 and X72) xor (X10 and X60 and X73) xor (X10 and X62 and X70) xor (X10 and X62 and X72) xor (X10 and X62 and X73) xor (X10 and X63 and X70) xor (X10 and X63 and X72) xor (X12 and X60 and X72) xor (X12 and X60 and X73) xor (X12 and X63 and X70) xor (X12 and X63 and X73) xor (X13 and X60 and X70) xor (X13 and X60 and X72) xor (X13 and X60 and X73) xor (X13 and X62 and X70) xor (X13 and X62 and X72) xor (X13 and X63 and X72) xor (X20 and X60 and X73) xor (X20 and X62 and X70) xor (X20 and X62 and X72) xor (X20 and X62 and X73) xor (X20 and X63 and X70) xor (X20 and X63 and X72) xor (X22 and X60 and X72) xor (X22 and X60 and X73) xor (X22 and X63 and X70) xor (X22 and X63 and X73) xor (X23 and X60 and X70) xor (X23 and X60 and X72) xor (X23 and X60 and X73) xor (X23 and X62 and X70) xor (X23 and X62 and X72) xor (X23 and X63 and X72) xor (X30 and X60 and X73) xor (X30 and X62 and X70) xor (X30 and X62 and X72) xor (X30 and X62 and X73) xor (X30 and X63 and X70) xor (X30 and X63 and X72) xor (X32 and X60 and X72) xor (X32 and X60 and X73) xor (X32 and X63 and X70) xor (X32 and X63 and X73) xor (X33 and X60 and X70) xor (X33 and X60 and X72) xor (X33 and X60 and X73) xor (X33 and X62 and X70) xor (X33 and X62 and X72) xor (X33 and X63 and X72) xor (X40 and X60 and X73) xor (X40 and X62 and X70) xor (X40 and X62 and X72) xor (X40 and X62 and X73) xor (X40 and X63 and X70) xor (X40 and X63 and X72) xor (X42 and X60 and X72) xor (X42 and X60 and X73) xor (X42 and X63 and X70) xor (X42 and X63 and X73) xor (X43 and X60 and X70) xor (X43 and X60 and X72) xor (X43 and X60 and X73) xor (X43 and X62 and X70) xor (X43 and X62 and X72) xor (X43 and X63 and X72) xor (X50 and X60 and X73) xor (X50 and X62 and X70) xor (X50 and X62 and X72) xor (X50 and X62 and X73) xor (X50 and X63 and X70) xor (X50 and X63 and X72) xor (X52 and X60 and X72) xor (X52 and X60 and X73) xor (X52 and X63 and X70) xor (X52 and X63 and X73) xor (X53 and X60 and X70) xor (X53 and X60 and X72) xor (X53 and X60 and X73) xor (X53 and X62 and X70) xor (X53 and X62 and X72) xor (X53 and X63 and X72));
    F53  <= ((X03 and X13) xor (X03 and X10) xor (X03 and X11) xor (X0_1 and X10) xor (X23) xor (X03 and X23) xor (X03 and X20) xor (X03 and X21) xor (X0_1 and X20) xor (X03 and X33) xor (X03 and X30) xor (X03 and X31) xor (X0_1 and X30) xor (X00 and X10 and X31) xor (X00 and X11 and X30) xor (X00 and X11 and X33) xor (X00 and X13 and X31) xor (X00 and X13 and X33) xor (X0_1 and X10 and X31) xor (X0_1 and X10 and X33) xor (X0_1 and X11 and X33) xor (X0_1 and X13 and X30) xor (X0_1 and X13 and X31) xor (X0_1 and X13 and X33) xor (X03 and X10 and X31) xor (X03 and X11 and X30) xor (X03 and X11 and X31) xor (X03 and X11 and X33) xor (X03 and X13 and X30) xor (X03 and X43) xor (X03 and X40) xor (X03 and X41) xor (X0_1 and X40) xor (X23 and X43) xor (X23 and X40) xor (X23 and X41) xor (X21 and X40) xor (X00 and X20 and X41) xor (X00 and X21 and X40) xor (X00 and X21 and X43) xor (X00 and X23 and X41) xor (X00 and X23 and X43) xor (X0_1 and X20 and X41) xor (X0_1 and X20 and X43) xor (X0_1 and X21 and X43) xor (X0_1 and X23 and X40) xor (X0_1 and X23 and X41) xor (X0_1 and X23 and X43) xor (X03 and X20 and X41) xor (X03 and X21 and X40) xor (X03 and X21 and X41) xor (X03 and X21 and X43) xor (X03 and X23 and X40) xor (X10 and X20 and X41) xor (X10 and X21 and X40) xor (X10 and X21 and X43) xor (X10 and X23 and X41) xor (X10 and X23 and X43) xor (X11 and X20 and X41) xor (X11 and X20 and X43) xor (X11 and X21 and X43) xor (X11 and X23 and X40) xor (X11 and X23 and X41) xor (X11 and X23 and X43) xor (X13 and X20 and X41) xor (X13 and X21 and X40) xor (X13 and X21 and X41) xor (X13 and X21 and X43) xor (X13 and X23 and X40) xor (X33 and X43) xor (X33 and X40) xor (X33 and X41) xor (X31 and X40) xor (X53) xor (X03 and X53) xor (X03 and X50) xor (X03 and X51) xor (X0_1 and X50) xor (X00 and X10 and X51) xor (X00 and X11 and X50) xor (X00 and X11 and X53) xor (X00 and X13 and X51) xor (X00 and X13 and X53) xor (X0_1 and X10 and X51) xor (X0_1 and X10 and X53) xor (X0_1 and X11 and X53) xor (X0_1 and X13 and X50) xor (X0_1 and X13 and X51) xor (X0_1 and X13 and X53) xor (X03 and X10 and X51) xor (X03 and X11 and X50) xor (X03 and X11 and X51) xor (X03 and X11 and X53) xor (X03 and X13 and X50) xor (X23 and X53) xor (X23 and X50) xor (X23 and X51) xor (X21 and X50) xor (X33 and X53) xor (X33 and X50) xor (X33 and X51) xor (X31 and X50) xor (X10 and X30 and X51) xor (X10 and X31 and X50) xor (X10 and X31 and X53) xor (X10 and X33 and X51) xor (X10 and X33 and X53) xor (X11 and X30 and X51) xor (X11 and X30 and X53) xor (X11 and X31 and X53) xor (X11 and X33 and X50) xor (X11 and X33 and X51) xor (X11 and X33 and X53) xor (X13 and X30 and X51) xor (X13 and X31 and X50) xor (X13 and X31 and X51) xor (X13 and X31 and X53) xor (X13 and X33 and X50) xor (X43 and X53) xor (X43 and X50) xor (X43 and X51) xor (X41 and X50) xor (X13 and X63) xor (X13 and X60) xor (X13 and X61) xor (X11 and X60) xor (X00 and X20 and X61) xor (X00 and X21 and X60) xor (X00 and X21 and X63) xor (X00 and X23 and X61) xor (X00 and X23 and X63) xor (X0_1 and X20 and X61) xor (X0_1 and X20 and X63) xor (X0_1 and X21 and X63) xor (X0_1 and X23 and X60) xor (X0_1 and X23 and X61) xor (X0_1 and X23 and X63) xor (X03 and X20 and X61) xor (X03 and X21 and X60) xor (X03 and X21 and X61) xor (X03 and X21 and X63) xor (X03 and X23 and X60) xor (X33 and X63) xor (X33 and X60) xor (X33 and X61) xor (X31 and X60) xor (X10 and X30 and X61) xor (X10 and X31 and X60) xor (X10 and X31 and X63) xor (X10 and X33 and X61) xor (X10 and X33 and X63) xor (X11 and X30 and X61) xor (X11 and X30 and X63) xor (X11 and X31 and X63) xor (X11 and X33 and X60) xor (X11 and X33 and X61) xor (X11 and X33 and X63) xor (X13 and X30 and X61) xor (X13 and X31 and X60) xor (X13 and X31 and X61) xor (X13 and X31 and X63) xor (X13 and X33 and X60) xor (X43 and X63) xor (X43 and X60) xor (X43 and X61) xor (X41 and X60) xor (X00 and X40 and X61) xor (X00 and X41 and X60) xor (X00 and X41 and X63) xor (X00 and X43 and X61) xor (X00 and X43 and X63) xor (X0_1 and X40 and X61) xor (X0_1 and X40 and X63) xor (X0_1 and X41 and X63) xor (X0_1 and X43 and X60) xor (X0_1 and X43 and X61) xor (X0_1 and X43 and X63) xor (X03 and X40 and X61) xor (X03 and X41 and X60) xor (X03 and X41 and X61) xor (X03 and X41 and X63) xor (X03 and X43 and X60) xor (X10 and X40 and X61) xor (X10 and X41 and X60) xor (X10 and X41 and X63) xor (X10 and X43 and X61) xor (X10 and X43 and X63) xor (X11 and X40 and X61) xor (X11 and X40 and X63) xor (X11 and X41 and X63) xor (X11 and X43 and X60) xor (X11 and X43 and X61) xor (X11 and X43 and X63) xor (X13 and X40 and X61) xor (X13 and X41 and X60) xor (X13 and X41 and X61) xor (X13 and X41 and X63) xor (X13 and X43 and X60) xor (X20 and X40 and X61) xor (X20 and X41 and X60) xor (X20 and X41 and X63) xor (X20 and X43 and X61) xor (X20 and X43 and X63) xor (X21 and X40 and X61) xor (X21 and X40 and X63) xor (X21 and X41 and X63) xor (X21 and X43 and X60) xor (X21 and X43 and X61) xor (X21 and X43 and X63) xor (X23 and X40 and X61) xor (X23 and X41 and X60) xor (X23 and X41 and X61) xor (X23 and X41 and X63) xor (X23 and X43 and X60) xor (X53 and X63) xor (X53 and X60) xor (X53 and X61) xor (X51 and X60) xor (X10 and X50 and X61) xor (X10 and X51 and X60) xor (X10 and X51 and X63) xor (X10 and X53 and X61) xor (X10 and X53 and X63) xor (X11 and X50 and X61) xor (X11 and X50 and X63) xor (X11 and X51 and X63) xor (X11 and X53 and X60) xor (X11 and X53 and X61) xor (X11 and X53 and X63) xor (X13 and X50 and X61) xor (X13 and X51 and X60) xor (X13 and X51 and X61) xor (X13 and X51 and X63) xor (X13 and X53 and X60) xor (X20 and X50 and X61) xor (X20 and X51 and X60) xor (X20 and X51 and X63) xor (X20 and X53 and X61) xor (X20 and X53 and X63) xor (X21 and X50 and X61) xor (X21 and X50 and X63) xor (X21 and X51 and X63) xor (X21 and X53 and X60) xor (X21 and X53 and X61) xor (X21 and X53 and X63) xor (X23 and X50 and X61) xor (X23 and X51 and X60) xor (X23 and X51 and X61) xor (X23 and X51 and X63) xor (X23 and X53 and X60) xor (X40 and X50 and X61) xor (X40 and X51 and X60) xor (X40 and X51 and X63) xor (X40 and X53 and X61) xor (X40 and X53 and X63) xor (X41 and X50 and X61) xor (X41 and X50 and X63) xor (X41 and X51 and X63) xor (X41 and X53 and X60) xor (X41 and X53 and X61) xor (X41 and X53 and X63) xor (X43 and X50 and X61) xor (X43 and X51 and X60) xor (X43 and X51 and X61) xor (X43 and X51 and X63) xor (X43 and X53 and X60) xor (X13 and X73) xor (X13 and X70) xor (X13 and X71) xor (X11 and X70) xor (X23 and X73) xor (X23 and X70) xor (X23 and X71) xor (X21 and X70) xor (X33 and X73) xor (X33 and X70) xor (X33 and X71) xor (X31 and X70) xor (X00 and X30 and X71) xor (X00 and X31 and X70) xor (X00 and X31 and X73) xor (X00 and X33 and X71) xor (X00 and X33 and X73) xor (X0_1 and X30 and X71) xor (X0_1 and X30 and X73) xor (X0_1 and X31 and X73) xor (X0_1 and X33 and X70) xor (X0_1 and X33 and X71) xor (X0_1 and X33 and X73) xor (X03 and X30 and X71) xor (X03 and X31 and X70) xor (X03 and X31 and X71) xor (X03 and X31 and X73) xor (X03 and X33 and X70) xor (X10 and X30 and X71) xor (X10 and X31 and X70) xor (X10 and X31 and X73) xor (X10 and X33 and X71) xor (X10 and X33 and X73) xor (X11 and X30 and X71) xor (X11 and X30 and X73) xor (X11 and X31 and X73) xor (X11 and X33 and X70) xor (X11 and X33 and X71) xor (X11 and X33 and X73) xor (X13 and X30 and X71) xor (X13 and X31 and X70) xor (X13 and X31 and X71) xor (X13 and X31 and X73) xor (X13 and X33 and X70) xor (X00 and X40 and X71) xor (X00 and X41 and X70) xor (X00 and X41 and X73) xor (X00 and X43 and X71) xor (X00 and X43 and X73) xor (X0_1 and X40 and X71) xor (X0_1 and X40 and X73) xor (X0_1 and X41 and X73) xor (X0_1 and X43 and X70) xor (X0_1 and X43 and X71) xor (X0_1 and X43 and X73) xor (X03 and X40 and X71) xor (X03 and X41 and X70) xor (X03 and X41 and X71) xor (X03 and X41 and X73) xor (X03 and X43 and X70) xor (X00 and X50 and X71) xor (X00 and X51 and X70) xor (X00 and X51 and X73) xor (X00 and X53 and X71) xor (X00 and X53 and X73) xor (X0_1 and X50 and X71) xor (X0_1 and X50 and X73) xor (X0_1 and X51 and X73) xor (X0_1 and X53 and X70) xor (X0_1 and X53 and X71) xor (X0_1 and X53 and X73) xor (X03 and X50 and X71) xor (X03 and X51 and X70) xor (X03 and X51 and X71) xor (X03 and X51 and X73) xor (X03 and X53 and X70) xor (X10 and X50 and X71) xor (X10 and X51 and X70) xor (X10 and X51 and X73) xor (X10 and X53 and X71) xor (X10 and X53 and X73) xor (X11 and X50 and X71) xor (X11 and X50 and X73) xor (X11 and X51 and X73) xor (X11 and X53 and X70) xor (X11 and X53 and X71) xor (X11 and X53 and X73) xor (X13 and X50 and X71) xor (X13 and X51 and X70) xor (X13 and X51 and X71) xor (X13 and X51 and X73) xor (X13 and X53 and X70) xor (X20 and X50 and X71) xor (X20 and X51 and X70) xor (X20 and X51 and X73) xor (X20 and X53 and X71) xor (X20 and X53 and X73) xor (X21 and X50 and X71) xor (X21 and X50 and X73) xor (X21 and X51 and X73) xor (X21 and X53 and X70) xor (X21 and X53 and X71) xor (X21 and X53 and X73) xor (X23 and X50 and X71) xor (X23 and X51 and X70) xor (X23 and X51 and X71) xor (X23 and X51 and X73) xor (X23 and X53 and X70) xor (X30 and X50 and X71) xor (X30 and X51 and X70) xor (X30 and X51 and X73) xor (X30 and X53 and X71) xor (X30 and X53 and X73) xor (X31 and X50 and X71) xor (X31 and X50 and X73) xor (X31 and X51 and X73) xor (X31 and X53 and X70) xor (X31 and X53 and X71) xor (X31 and X53 and X73) xor (X33 and X50 and X71) xor (X33 and X51 and X70) xor (X33 and X51 and X71) xor (X33 and X51 and X73) xor (X33 and X53 and X70) xor (X10 and X60 and X71) xor (X10 and X61 and X70) xor (X10 and X61 and X73) xor (X10 and X63 and X71) xor (X10 and X63 and X73) xor (X11 and X60 and X71) xor (X11 and X60 and X73) xor (X11 and X61 and X73) xor (X11 and X63 and X70) xor (X11 and X63 and X71) xor (X11 and X63 and X73) xor (X13 and X60 and X71) xor (X13 and X61 and X70) xor (X13 and X61 and X71) xor (X13 and X61 and X73) xor (X13 and X63 and X70) xor (X20 and X60 and X71) xor (X20 and X61 and X70) xor (X20 and X61 and X73) xor (X20 and X63 and X71) xor (X20 and X63 and X73) xor (X21 and X60 and X71) xor (X21 and X60 and X73) xor (X21 and X61 and X73) xor (X21 and X63 and X70) xor (X21 and X63 and X71) xor (X21 and X63 and X73) xor (X23 and X60 and X71) xor (X23 and X61 and X70) xor (X23 and X61 and X71) xor (X23 and X61 and X73) xor (X23 and X63 and X70) xor (X30 and X60 and X71) xor (X30 and X61 and X70) xor (X30 and X61 and X73) xor (X30 and X63 and X71) xor (X30 and X63 and X73) xor (X31 and X60 and X71) xor (X31 and X60 and X73) xor (X31 and X61 and X73) xor (X31 and X63 and X70) xor (X31 and X63 and X71) xor (X31 and X63 and X73) xor (X33 and X60 and X71) xor (X33 and X61 and X70) xor (X33 and X61 and X71) xor (X33 and X61 and X73) xor (X33 and X63 and X70) xor (X40 and X60 and X71) xor (X40 and X61 and X70) xor (X40 and X61 and X73) xor (X40 and X63 and X71) xor (X40 and X63 and X73) xor (X41 and X60 and X71) xor (X41 and X60 and X73) xor (X41 and X61 and X73) xor (X41 and X63 and X70) xor (X41 and X63 and X71) xor (X41 and X63 and X73) xor (X43 and X60 and X71) xor (X43 and X61 and X70) xor (X43 and X61 and X71) xor (X43 and X61 and X73) xor (X43 and X63 and X70) xor (X50 and X60 and X71) xor (X50 and X61 and X70) xor (X50 and X61 and X73) xor (X50 and X63 and X71) xor (X50 and X63 and X73) xor (X51 and X60 and X71) xor (X51 and X60 and X73) xor (X51 and X61 and X73) xor (X51 and X63 and X70) xor (X51 and X63 and X71) xor (X51 and X63 and X73) xor (X53 and X60 and X71) xor (X53 and X61 and X70) xor (X53 and X61 and X71) xor (X53 and X61 and X73) xor (X53 and X63 and X70));
    F60  <= ((X10) xor (X20) xor (X10 and X20) xor (X10 and X21) xor (X12 and X20) xor (X10 and X22) xor (X00 and X10 and X20) xor (X00 and X10 and X22) xor (X00 and X11 and X21) xor (X00 and X11 and X22) xor (X00 and X12 and X21) xor (X0_1 and X10 and X20) xor (X0_1 and X10 and X22) xor (X0_1 and X11 and X20) xor (X0_1 and X12 and X20) xor (X0_1 and X12 and X21) xor (X02 and X10 and X20) xor (X02 and X10 and X21) xor (X02 and X11 and X20) xor (X02 and X11 and X21) xor (X02 and X12 and X20) xor (X02 and X12 and X22) xor (X00 and X30) xor (X00 and X31) xor (X02 and X30) xor (X00 and X32) xor (X20 and X30) xor (X20 and X31) xor (X22 and X30) xor (X20 and X32) xor (X00 and X20 and X30) xor (X00 and X20 and X32) xor (X00 and X21 and X31) xor (X00 and X21 and X32) xor (X00 and X22 and X31) xor (X0_1 and X20 and X30) xor (X0_1 and X20 and X32) xor (X0_1 and X21 and X30) xor (X0_1 and X22 and X30) xor (X0_1 and X22 and X31) xor (X02 and X20 and X30) xor (X02 and X20 and X31) xor (X02 and X21 and X30) xor (X02 and X21 and X31) xor (X02 and X22 and X30) xor (X02 and X22 and X32) xor (X10 and X20 and X30) xor (X10 and X20 and X32) xor (X10 and X21 and X31) xor (X10 and X21 and X32) xor (X10 and X22 and X31) xor (X11 and X20 and X30) xor (X11 and X20 and X32) xor (X11 and X21 and X30) xor (X11 and X22 and X30) xor (X11 and X22 and X31) xor (X12 and X20 and X30) xor (X12 and X20 and X31) xor (X12 and X21 and X30) xor (X12 and X21 and X31) xor (X12 and X22 and X30) xor (X12 and X22 and X32) xor (X40) xor (X00 and X40) xor (X00 and X41) xor (X02 and X40) xor (X00 and X42) xor (X00 and X10 and X40) xor (X00 and X10 and X42) xor (X00 and X11 and X41) xor (X00 and X11 and X42) xor (X00 and X12 and X41) xor (X0_1 and X10 and X40) xor (X0_1 and X10 and X42) xor (X0_1 and X11 and X40) xor (X0_1 and X12 and X40) xor (X0_1 and X12 and X41) xor (X02 and X10 and X40) xor (X02 and X10 and X41) xor (X02 and X11 and X40) xor (X02 and X11 and X41) xor (X02 and X12 and X40) xor (X02 and X12 and X42) xor (X20 and X40) xor (X20 and X41) xor (X22 and X40) xor (X20 and X42) xor (X00 and X20 and X40) xor (X00 and X20 and X42) xor (X00 and X21 and X41) xor (X00 and X21 and X42) xor (X00 and X22 and X41) xor (X0_1 and X20 and X40) xor (X0_1 and X20 and X42) xor (X0_1 and X21 and X40) xor (X0_1 and X22 and X40) xor (X0_1 and X22 and X41) xor (X02 and X20 and X40) xor (X02 and X20 and X41) xor (X02 and X21 and X40) xor (X02 and X21 and X41) xor (X02 and X22 and X40) xor (X02 and X22 and X42) xor (X10 and X20 and X40) xor (X10 and X20 and X42) xor (X10 and X21 and X41) xor (X10 and X21 and X42) xor (X10 and X22 and X41) xor (X11 and X20 and X40) xor (X11 and X20 and X42) xor (X11 and X21 and X40) xor (X11 and X22 and X40) xor (X11 and X22 and X41) xor (X12 and X20 and X40) xor (X12 and X20 and X41) xor (X12 and X21 and X40) xor (X12 and X21 and X41) xor (X12 and X22 and X40) xor (X12 and X22 and X42) xor (X30 and X40) xor (X30 and X41) xor (X32 and X40) xor (X30 and X42) xor (X00 and X30 and X40) xor (X00 and X30 and X42) xor (X00 and X31 and X41) xor (X00 and X31 and X42) xor (X00 and X32 and X41) xor (X0_1 and X30 and X40) xor (X0_1 and X30 and X42) xor (X0_1 and X31 and X40) xor (X0_1 and X32 and X40) xor (X0_1 and X32 and X41) xor (X02 and X30 and X40) xor (X02 and X30 and X41) xor (X02 and X31 and X40) xor (X02 and X31 and X41) xor (X02 and X32 and X40) xor (X02 and X32 and X42) xor (X00 and X50) xor (X00 and X51) xor (X02 and X50) xor (X00 and X52) xor (X20 and X50) xor (X20 and X51) xor (X22 and X50) xor (X20 and X52) xor (X10 and X20 and X50) xor (X10 and X20 and X52) xor (X10 and X21 and X51) xor (X10 and X21 and X52) xor (X10 and X22 and X51) xor (X11 and X20 and X50) xor (X11 and X20 and X52) xor (X11 and X21 and X50) xor (X11 and X22 and X50) xor (X11 and X22 and X51) xor (X12 and X20 and X50) xor (X12 and X20 and X51) xor (X12 and X21 and X50) xor (X12 and X21 and X51) xor (X12 and X22 and X50) xor (X12 and X22 and X52) xor (X00 and X30 and X50) xor (X00 and X30 and X52) xor (X00 and X31 and X51) xor (X00 and X31 and X52) xor (X00 and X32 and X51) xor (X0_1 and X30 and X50) xor (X0_1 and X30 and X52) xor (X0_1 and X31 and X50) xor (X0_1 and X32 and X50) xor (X0_1 and X32 and X51) xor (X02 and X30 and X50) xor (X02 and X30 and X51) xor (X02 and X31 and X50) xor (X02 and X31 and X51) xor (X02 and X32 and X50) xor (X02 and X32 and X52) xor (X40 and X50) xor (X40 and X51) xor (X42 and X50) xor (X40 and X52) xor (X30 and X40 and X50) xor (X30 and X40 and X52) xor (X30 and X41 and X51) xor (X30 and X41 and X52) xor (X30 and X42 and X51) xor (X31 and X40 and X50) xor (X31 and X40 and X52) xor (X31 and X41 and X50) xor (X31 and X42 and X50) xor (X31 and X42 and X51) xor (X32 and X40 and X50) xor (X32 and X40 and X51) xor (X32 and X41 and X50) xor (X32 and X41 and X51) xor (X32 and X42 and X50) xor (X32 and X42 and X52) xor (X60) xor (X00 and X60) xor (X00 and X61) xor (X02 and X60) xor (X00 and X62) xor (X10 and X60) xor (X10 and X61) xor (X12 and X60) xor (X10 and X62) xor (X30 and X60) xor (X30 and X61) xor (X32 and X60) xor (X30 and X62) xor (X40 and X60) xor (X40 and X61) xor (X42 and X60) xor (X40 and X62) xor (X10 and X40 and X60) xor (X10 and X40 and X62) xor (X10 and X41 and X61) xor (X10 and X41 and X62) xor (X10 and X42 and X61) xor (X11 and X40 and X60) xor (X11 and X40 and X62) xor (X11 and X41 and X60) xor (X11 and X42 and X60) xor (X11 and X42 and X61) xor (X12 and X40 and X60) xor (X12 and X40 and X61) xor (X12 and X41 and X60) xor (X12 and X41 and X61) xor (X12 and X42 and X60) xor (X12 and X42 and X62) xor (X30 and X40 and X60) xor (X30 and X40 and X62) xor (X30 and X41 and X61) xor (X30 and X41 and X62) xor (X30 and X42 and X61) xor (X31 and X40 and X60) xor (X31 and X40 and X62) xor (X31 and X41 and X60) xor (X31 and X42 and X60) xor (X31 and X42 and X61) xor (X32 and X40 and X60) xor (X32 and X40 and X61) xor (X32 and X41 and X60) xor (X32 and X41 and X61) xor (X32 and X42 and X60) xor (X32 and X42 and X62) xor (X10 and X50 and X60) xor (X10 and X50 and X62) xor (X10 and X51 and X61) xor (X10 and X51 and X62) xor (X10 and X52 and X61) xor (X11 and X50 and X60) xor (X11 and X50 and X62) xor (X11 and X51 and X60) xor (X11 and X52 and X60) xor (X11 and X52 and X61) xor (X12 and X50 and X60) xor (X12 and X50 and X61) xor (X12 and X51 and X60) xor (X12 and X51 and X61) xor (X12 and X52 and X60) xor (X12 and X52 and X62) xor (X20 and X50 and X60) xor (X20 and X50 and X62) xor (X20 and X51 and X61) xor (X20 and X51 and X62) xor (X20 and X52 and X61) xor (X21 and X50 and X60) xor (X21 and X50 and X62) xor (X21 and X51 and X60) xor (X21 and X52 and X60) xor (X21 and X52 and X61) xor (X22 and X50 and X60) xor (X22 and X50 and X61) xor (X22 and X51 and X60) xor (X22 and X51 and X61) xor (X22 and X52 and X60) xor (X22 and X52 and X62) xor (X30 and X50 and X60) xor (X30 and X50 and X62) xor (X30 and X51 and X61) xor (X30 and X51 and X62) xor (X30 and X52 and X61) xor (X31 and X50 and X60) xor (X31 and X50 and X62) xor (X31 and X51 and X60) xor (X31 and X52 and X60) xor (X31 and X52 and X61) xor (X32 and X50 and X60) xor (X32 and X50 and X61) xor (X32 and X51 and X60) xor (X32 and X51 and X61) xor (X32 and X52 and X60) xor (X32 and X52 and X62) xor (X00 and X10 and X70) xor (X00 and X10 and X72) xor (X00 and X11 and X71) xor (X00 and X11 and X72) xor (X00 and X12 and X71) xor (X0_1 and X10 and X70) xor (X0_1 and X10 and X72) xor (X0_1 and X11 and X70) xor (X0_1 and X12 and X70) xor (X0_1 and X12 and X71) xor (X02 and X10 and X70) xor (X02 and X10 and X71) xor (X02 and X11 and X70) xor (X02 and X11 and X71) xor (X02 and X12 and X70) xor (X02 and X12 and X72) xor (X00 and X20 and X70) xor (X00 and X20 and X72) xor (X00 and X21 and X71) xor (X00 and X21 and X72) xor (X00 and X22 and X71) xor (X0_1 and X20 and X70) xor (X0_1 and X20 and X72) xor (X0_1 and X21 and X70) xor (X0_1 and X22 and X70) xor (X0_1 and X22 and X71) xor (X02 and X20 and X70) xor (X02 and X20 and X71) xor (X02 and X21 and X70) xor (X02 and X21 and X71) xor (X02 and X22 and X70) xor (X02 and X22 and X72) xor (X10 and X20 and X70) xor (X10 and X20 and X72) xor (X10 and X21 and X71) xor (X10 and X21 and X72) xor (X10 and X22 and X71) xor (X11 and X20 and X70) xor (X11 and X20 and X72) xor (X11 and X21 and X70) xor (X11 and X22 and X70) xor (X11 and X22 and X71) xor (X12 and X20 and X70) xor (X12 and X20 and X71) xor (X12 and X21 and X70) xor (X12 and X21 and X71) xor (X12 and X22 and X70) xor (X12 and X22 and X72) xor (X30 and X70) xor (X30 and X71) xor (X32 and X70) xor (X30 and X72) xor (X10 and X30 and X70) xor (X10 and X30 and X72) xor (X10 and X31 and X71) xor (X10 and X31 and X72) xor (X10 and X32 and X71) xor (X11 and X30 and X70) xor (X11 and X30 and X72) xor (X11 and X31 and X70) xor (X11 and X32 and X70) xor (X11 and X32 and X71) xor (X12 and X30 and X70) xor (X12 and X30 and X71) xor (X12 and X31 and X70) xor (X12 and X31 and X71) xor (X12 and X32 and X70) xor (X12 and X32 and X72) xor (X40 and X70) xor (X40 and X71) xor (X42 and X70) xor (X40 and X72) xor (X00 and X40 and X70) xor (X00 and X40 and X72) xor (X00 and X41 and X71) xor (X00 and X41 and X72) xor (X00 and X42 and X71) xor (X0_1 and X40 and X70) xor (X0_1 and X40 and X72) xor (X0_1 and X41 and X70) xor (X0_1 and X42 and X70) xor (X0_1 and X42 and X71) xor (X02 and X40 and X70) xor (X02 and X40 and X71) xor (X02 and X41 and X70) xor (X02 and X41 and X71) xor (X02 and X42 and X70) xor (X02 and X42 and X72) xor (X10 and X40 and X70) xor (X10 and X40 and X72) xor (X10 and X41 and X71) xor (X10 and X41 and X72) xor (X10 and X42 and X71) xor (X11 and X40 and X70) xor (X11 and X40 and X72) xor (X11 and X41 and X70) xor (X11 and X42 and X70) xor (X11 and X42 and X71) xor (X12 and X40 and X70) xor (X12 and X40 and X71) xor (X12 and X41 and X70) xor (X12 and X41 and X71) xor (X12 and X42 and X70) xor (X12 and X42 and X72) xor (X20 and X40 and X70) xor (X20 and X40 and X72) xor (X20 and X41 and X71) xor (X20 and X41 and X72) xor (X20 and X42 and X71) xor (X21 and X40 and X70) xor (X21 and X40 and X72) xor (X21 and X41 and X70) xor (X21 and X42 and X70) xor (X21 and X42 and X71) xor (X22 and X40 and X70) xor (X22 and X40 and X71) xor (X22 and X41 and X70) xor (X22 and X41 and X71) xor (X22 and X42 and X70) xor (X22 and X42 and X72) xor (X50 and X70) xor (X50 and X71) xor (X52 and X70) xor (X50 and X72) xor (X00 and X50 and X70) xor (X00 and X50 and X72) xor (X00 and X51 and X71) xor (X00 and X51 and X72) xor (X00 and X52 and X71) xor (X0_1 and X50 and X70) xor (X0_1 and X50 and X72) xor (X0_1 and X51 and X70) xor (X0_1 and X52 and X70) xor (X0_1 and X52 and X71) xor (X02 and X50 and X70) xor (X02 and X50 and X71) xor (X02 and X51 and X70) xor (X02 and X51 and X71) xor (X02 and X52 and X70) xor (X02 and X52 and X72) xor (X60 and X70) xor (X60 and X71) xor (X62 and X70) xor (X60 and X72) xor (X00 and X60 and X70) xor (X00 and X60 and X72) xor (X00 and X61 and X71) xor (X00 and X61 and X72) xor (X00 and X62 and X71) xor (X0_1 and X60 and X70) xor (X0_1 and X60 and X72) xor (X0_1 and X61 and X70) xor (X0_1 and X62 and X70) xor (X0_1 and X62 and X71) xor (X02 and X60 and X70) xor (X02 and X60 and X71) xor (X02 and X61 and X70) xor (X02 and X61 and X71) xor (X02 and X62 and X70) xor (X02 and X62 and X72) xor (X30 and X60 and X70) xor (X30 and X60 and X72) xor (X30 and X61 and X71) xor (X30 and X61 and X72) xor (X30 and X62 and X71) xor (X31 and X60 and X70) xor (X31 and X60 and X72) xor (X31 and X61 and X70) xor (X31 and X62 and X70) xor (X31 and X62 and X71) xor (X32 and X60 and X70) xor (X32 and X60 and X71) xor (X32 and X61 and X70) xor (X32 and X61 and X71) xor (X32 and X62 and X70) xor (X32 and X62 and X72));
    F61  <= ((X11) xor (X21) xor (X11 and X21) xor (X11 and X22) xor (X12 and X21) xor (X11 and X23) xor (X0_1 and X11 and X21) xor (X0_1 and X11 and X22) xor (X0_1 and X12 and X22) xor (X0_1 and X12 and X23) xor (X0_1 and X13 and X22) xor (X02 and X11 and X22) xor (X02 and X11 and X23) xor (X02 and X12 and X21) xor (X02 and X12 and X23) xor (X02 and X13 and X21) xor (X02 and X13 and X22) xor (X03 and X11 and X22) xor (X03 and X12 and X21) xor (X03 and X12 and X23) xor (X03 and X13 and X21) xor (X03 and X13 and X23) xor (X0_1 and X31) xor (X0_1 and X32) xor (X02 and X31) xor (X0_1 and X33) xor (X21 and X31) xor (X21 and X32) xor (X22 and X31) xor (X21 and X33) xor (X0_1 and X21 and X31) xor (X0_1 and X21 and X32) xor (X0_1 and X22 and X32) xor (X0_1 and X22 and X33) xor (X0_1 and X23 and X32) xor (X02 and X21 and X32) xor (X02 and X21 and X33) xor (X02 and X22 and X31) xor (X02 and X22 and X33) xor (X02 and X23 and X31) xor (X02 and X23 and X32) xor (X03 and X21 and X32) xor (X03 and X22 and X31) xor (X03 and X22 and X33) xor (X03 and X23 and X31) xor (X03 and X23 and X33) xor (X11 and X21 and X31) xor (X11 and X21 and X32) xor (X11 and X22 and X32) xor (X11 and X22 and X33) xor (X11 and X23 and X32) xor (X12 and X21 and X32) xor (X12 and X21 and X33) xor (X12 and X22 and X31) xor (X12 and X22 and X33) xor (X12 and X23 and X31) xor (X12 and X23 and X32) xor (X13 and X21 and X32) xor (X13 and X22 and X31) xor (X13 and X22 and X33) xor (X13 and X23 and X31) xor (X13 and X23 and X33) xor (X41) xor (X0_1 and X41) xor (X0_1 and X42) xor (X02 and X41) xor (X0_1 and X43) xor (X0_1 and X11 and X41) xor (X0_1 and X11 and X42) xor (X0_1 and X12 and X42) xor (X0_1 and X12 and X43) xor (X0_1 and X13 and X42) xor (X02 and X11 and X42) xor (X02 and X11 and X43) xor (X02 and X12 and X41) xor (X02 and X12 and X43) xor (X02 and X13 and X41) xor (X02 and X13 and X42) xor (X03 and X11 and X42) xor (X03 and X12 and X41) xor (X03 and X12 and X43) xor (X03 and X13 and X41) xor (X03 and X13 and X43) xor (X21 and X41) xor (X21 and X42) xor (X22 and X41) xor (X21 and X43) xor (X0_1 and X21 and X41) xor (X0_1 and X21 and X42) xor (X0_1 and X22 and X42) xor (X0_1 and X22 and X43) xor (X0_1 and X23 and X42) xor (X02 and X21 and X42) xor (X02 and X21 and X43) xor (X02 and X22 and X41) xor (X02 and X22 and X43) xor (X02 and X23 and X41) xor (X02 and X23 and X42) xor (X03 and X21 and X42) xor (X03 and X22 and X41) xor (X03 and X22 and X43) xor (X03 and X23 and X41) xor (X03 and X23 and X43) xor (X11 and X21 and X41) xor (X11 and X21 and X42) xor (X11 and X22 and X42) xor (X11 and X22 and X43) xor (X11 and X23 and X42) xor (X12 and X21 and X42) xor (X12 and X21 and X43) xor (X12 and X22 and X41) xor (X12 and X22 and X43) xor (X12 and X23 and X41) xor (X12 and X23 and X42) xor (X13 and X21 and X42) xor (X13 and X22 and X41) xor (X13 and X22 and X43) xor (X13 and X23 and X41) xor (X13 and X23 and X43) xor (X31 and X41) xor (X31 and X42) xor (X32 and X41) xor (X31 and X43) xor (X0_1 and X31 and X41) xor (X0_1 and X31 and X42) xor (X0_1 and X32 and X42) xor (X0_1 and X32 and X43) xor (X0_1 and X33 and X42) xor (X02 and X31 and X42) xor (X02 and X31 and X43) xor (X02 and X32 and X41) xor (X02 and X32 and X43) xor (X02 and X33 and X41) xor (X02 and X33 and X42) xor (X03 and X31 and X42) xor (X03 and X32 and X41) xor (X03 and X32 and X43) xor (X03 and X33 and X41) xor (X03 and X33 and X43) xor (X0_1 and X51) xor (X0_1 and X52) xor (X02 and X51) xor (X0_1 and X53) xor (X21 and X51) xor (X21 and X52) xor (X22 and X51) xor (X21 and X53) xor (X11 and X21 and X51) xor (X11 and X21 and X52) xor (X11 and X22 and X52) xor (X11 and X22 and X53) xor (X11 and X23 and X52) xor (X12 and X21 and X52) xor (X12 and X21 and X53) xor (X12 and X22 and X51) xor (X12 and X22 and X53) xor (X12 and X23 and X51) xor (X12 and X23 and X52) xor (X13 and X21 and X52) xor (X13 and X22 and X51) xor (X13 and X22 and X53) xor (X13 and X23 and X51) xor (X13 and X23 and X53) xor (X0_1 and X31 and X51) xor (X0_1 and X31 and X52) xor (X0_1 and X32 and X52) xor (X0_1 and X32 and X53) xor (X0_1 and X33 and X52) xor (X02 and X31 and X52) xor (X02 and X31 and X53) xor (X02 and X32 and X51) xor (X02 and X32 and X53) xor (X02 and X33 and X51) xor (X02 and X33 and X52) xor (X03 and X31 and X52) xor (X03 and X32 and X51) xor (X03 and X32 and X53) xor (X03 and X33 and X51) xor (X03 and X33 and X53) xor (X41 and X51) xor (X41 and X52) xor (X42 and X51) xor (X41 and X53) xor (X31 and X41 and X51) xor (X31 and X41 and X52) xor (X31 and X42 and X52) xor (X31 and X42 and X53) xor (X31 and X43 and X52) xor (X32 and X41 and X52) xor (X32 and X41 and X53) xor (X32 and X42 and X51) xor (X32 and X42 and X53) xor (X32 and X43 and X51) xor (X32 and X43 and X52) xor (X33 and X41 and X52) xor (X33 and X42 and X51) xor (X33 and X42 and X53) xor (X33 and X43 and X51) xor (X33 and X43 and X53) xor (X61) xor (X0_1 and X61) xor (X0_1 and X62) xor (X02 and X61) xor (X0_1 and X63) xor (X11 and X61) xor (X11 and X62) xor (X12 and X61) xor (X11 and X63) xor (X31 and X61) xor (X31 and X62) xor (X32 and X61) xor (X31 and X63) xor (X41 and X61) xor (X41 and X62) xor (X42 and X61) xor (X41 and X63) xor (X11 and X41 and X61) xor (X11 and X41 and X62) xor (X11 and X42 and X62) xor (X11 and X42 and X63) xor (X11 and X43 and X62) xor (X12 and X41 and X62) xor (X12 and X41 and X63) xor (X12 and X42 and X61) xor (X12 and X42 and X63) xor (X12 and X43 and X61) xor (X12 and X43 and X62) xor (X13 and X41 and X62) xor (X13 and X42 and X61) xor (X13 and X42 and X63) xor (X13 and X43 and X61) xor (X13 and X43 and X63) xor (X31 and X41 and X61) xor (X31 and X41 and X62) xor (X31 and X42 and X62) xor (X31 and X42 and X63) xor (X31 and X43 and X62) xor (X32 and X41 and X62) xor (X32 and X41 and X63) xor (X32 and X42 and X61) xor (X32 and X42 and X63) xor (X32 and X43 and X61) xor (X32 and X43 and X62) xor (X33 and X41 and X62) xor (X33 and X42 and X61) xor (X33 and X42 and X63) xor (X33 and X43 and X61) xor (X33 and X43 and X63) xor (X11 and X51 and X61) xor (X11 and X51 and X62) xor (X11 and X52 and X62) xor (X11 and X52 and X63) xor (X11 and X53 and X62) xor (X12 and X51 and X62) xor (X12 and X51 and X63) xor (X12 and X52 and X61) xor (X12 and X52 and X63) xor (X12 and X53 and X61) xor (X12 and X53 and X62) xor (X13 and X51 and X62) xor (X13 and X52 and X61) xor (X13 and X52 and X63) xor (X13 and X53 and X61) xor (X13 and X53 and X63) xor (X21 and X51 and X61) xor (X21 and X51 and X62) xor (X21 and X52 and X62) xor (X21 and X52 and X63) xor (X21 and X53 and X62) xor (X22 and X51 and X62) xor (X22 and X51 and X63) xor (X22 and X52 and X61) xor (X22 and X52 and X63) xor (X22 and X53 and X61) xor (X22 and X53 and X62) xor (X23 and X51 and X62) xor (X23 and X52 and X61) xor (X23 and X52 and X63) xor (X23 and X53 and X61) xor (X23 and X53 and X63) xor (X31 and X51 and X61) xor (X31 and X51 and X62) xor (X31 and X52 and X62) xor (X31 and X52 and X63) xor (X31 and X53 and X62) xor (X32 and X51 and X62) xor (X32 and X51 and X63) xor (X32 and X52 and X61) xor (X32 and X52 and X63) xor (X32 and X53 and X61) xor (X32 and X53 and X62) xor (X33 and X51 and X62) xor (X33 and X52 and X61) xor (X33 and X52 and X63) xor (X33 and X53 and X61) xor (X33 and X53 and X63) xor (X0_1 and X11 and X71) xor (X0_1 and X11 and X72) xor (X0_1 and X12 and X72) xor (X0_1 and X12 and X73) xor (X0_1 and X13 and X72) xor (X02 and X11 and X72) xor (X02 and X11 and X73) xor (X02 and X12 and X71) xor (X02 and X12 and X73) xor (X02 and X13 and X71) xor (X02 and X13 and X72) xor (X03 and X11 and X72) xor (X03 and X12 and X71) xor (X03 and X12 and X73) xor (X03 and X13 and X71) xor (X03 and X13 and X73) xor (X0_1 and X21 and X71) xor (X0_1 and X21 and X72) xor (X0_1 and X22 and X72) xor (X0_1 and X22 and X73) xor (X0_1 and X23 and X72) xor (X02 and X21 and X72) xor (X02 and X21 and X73) xor (X02 and X22 and X71) xor (X02 and X22 and X73) xor (X02 and X23 and X71) xor (X02 and X23 and X72) xor (X03 and X21 and X72) xor (X03 and X22 and X71) xor (X03 and X22 and X73) xor (X03 and X23 and X71) xor (X03 and X23 and X73) xor (X11 and X21 and X71) xor (X11 and X21 and X72) xor (X11 and X22 and X72) xor (X11 and X22 and X73) xor (X11 and X23 and X72) xor (X12 and X21 and X72) xor (X12 and X21 and X73) xor (X12 and X22 and X71) xor (X12 and X22 and X73) xor (X12 and X23 and X71) xor (X12 and X23 and X72) xor (X13 and X21 and X72) xor (X13 and X22 and X71) xor (X13 and X22 and X73) xor (X13 and X23 and X71) xor (X13 and X23 and X73) xor (X31 and X71) xor (X31 and X72) xor (X32 and X71) xor (X31 and X73) xor (X11 and X31 and X71) xor (X11 and X31 and X72) xor (X11 and X32 and X72) xor (X11 and X32 and X73) xor (X11 and X33 and X72) xor (X12 and X31 and X72) xor (X12 and X31 and X73) xor (X12 and X32 and X71) xor (X12 and X32 and X73) xor (X12 and X33 and X71) xor (X12 and X33 and X72) xor (X13 and X31 and X72) xor (X13 and X32 and X71) xor (X13 and X32 and X73) xor (X13 and X33 and X71) xor (X13 and X33 and X73) xor (X41 and X71) xor (X41 and X72) xor (X42 and X71) xor (X41 and X73) xor (X0_1 and X41 and X71) xor (X0_1 and X41 and X72) xor (X0_1 and X42 and X72) xor (X0_1 and X42 and X73) xor (X0_1 and X43 and X72) xor (X02 and X41 and X72) xor (X02 and X41 and X73) xor (X02 and X42 and X71) xor (X02 and X42 and X73) xor (X02 and X43 and X71) xor (X02 and X43 and X72) xor (X03 and X41 and X72) xor (X03 and X42 and X71) xor (X03 and X42 and X73) xor (X03 and X43 and X71) xor (X03 and X43 and X73) xor (X11 and X41 and X71) xor (X11 and X41 and X72) xor (X11 and X42 and X72) xor (X11 and X42 and X73) xor (X11 and X43 and X72) xor (X12 and X41 and X72) xor (X12 and X41 and X73) xor (X12 and X42 and X71) xor (X12 and X42 and X73) xor (X12 and X43 and X71) xor (X12 and X43 and X72) xor (X13 and X41 and X72) xor (X13 and X42 and X71) xor (X13 and X42 and X73) xor (X13 and X43 and X71) xor (X13 and X43 and X73) xor (X21 and X41 and X71) xor (X21 and X41 and X72) xor (X21 and X42 and X72) xor (X21 and X42 and X73) xor (X21 and X43 and X72) xor (X22 and X41 and X72) xor (X22 and X41 and X73) xor (X22 and X42 and X71) xor (X22 and X42 and X73) xor (X22 and X43 and X71) xor (X22 and X43 and X72) xor (X23 and X41 and X72) xor (X23 and X42 and X71) xor (X23 and X42 and X73) xor (X23 and X43 and X71) xor (X23 and X43 and X73) xor (X51 and X71) xor (X51 and X72) xor (X52 and X71) xor (X51 and X73) xor (X0_1 and X51 and X71) xor (X0_1 and X51 and X72) xor (X0_1 and X52 and X72) xor (X0_1 and X52 and X73) xor (X0_1 and X53 and X72) xor (X02 and X51 and X72) xor (X02 and X51 and X73) xor (X02 and X52 and X71) xor (X02 and X52 and X73) xor (X02 and X53 and X71) xor (X02 and X53 and X72) xor (X03 and X51 and X72) xor (X03 and X52 and X71) xor (X03 and X52 and X73) xor (X03 and X53 and X71) xor (X03 and X53 and X73) xor (X61 and X71) xor (X61 and X72) xor (X62 and X71) xor (X61 and X73) xor (X0_1 and X61 and X71) xor (X0_1 and X61 and X72) xor (X0_1 and X62 and X72) xor (X0_1 and X62 and X73) xor (X0_1 and X63 and X72) xor (X02 and X61 and X72) xor (X02 and X61 and X73) xor (X02 and X62 and X71) xor (X02 and X62 and X73) xor (X02 and X63 and X71) xor (X02 and X63 and X72) xor (X03 and X61 and X72) xor (X03 and X62 and X71) xor (X03 and X62 and X73) xor (X03 and X63 and X71) xor (X03 and X63 and X73) xor (X31 and X61 and X71) xor (X31 and X61 and X72) xor (X31 and X62 and X72) xor (X31 and X62 and X73) xor (X31 and X63 and X72) xor (X32 and X61 and X72) xor (X32 and X61 and X73) xor (X32 and X62 and X71) xor (X32 and X62 and X73) xor (X32 and X63 and X71) xor (X32 and X63 and X72) xor (X33 and X61 and X72) xor (X33 and X62 and X71) xor (X33 and X62 and X73) xor (X33 and X63 and X71) xor (X33 and X63 and X73));
    F62  <= ((X12) xor (X22) xor (X12 and X22) xor (X10 and X23) xor (X12 and X23) xor (X13 and X22) xor (X00 and X10 and X23) xor (X00 and X12 and X20) xor (X00 and X12 and X22) xor (X00 and X12 and X23) xor (X00 and X13 and X20) xor (X00 and X13 and X22) xor (X02 and X10 and X22) xor (X02 and X10 and X23) xor (X02 and X13 and X20) xor (X02 and X13 and X23) xor (X03 and X10 and X20) xor (X03 and X10 and X22) xor (X03 and X10 and X23) xor (X03 and X12 and X20) xor (X03 and X12 and X22) xor (X03 and X13 and X22) xor (X02 and X32) xor (X00 and X33) xor (X02 and X33) xor (X03 and X32) xor (X22 and X32) xor (X20 and X33) xor (X22 and X33) xor (X23 and X32) xor (X00 and X20 and X33) xor (X00 and X22 and X30) xor (X00 and X22 and X32) xor (X00 and X22 and X33) xor (X00 and X23 and X30) xor (X00 and X23 and X32) xor (X02 and X20 and X32) xor (X02 and X20 and X33) xor (X02 and X23 and X30) xor (X02 and X23 and X33) xor (X03 and X20 and X30) xor (X03 and X20 and X32) xor (X03 and X20 and X33) xor (X03 and X22 and X30) xor (X03 and X22 and X32) xor (X03 and X23 and X32) xor (X10 and X20 and X33) xor (X10 and X22 and X30) xor (X10 and X22 and X32) xor (X10 and X22 and X33) xor (X10 and X23 and X30) xor (X10 and X23 and X32) xor (X12 and X20 and X32) xor (X12 and X20 and X33) xor (X12 and X23 and X30) xor (X12 and X23 and X33) xor (X13 and X20 and X30) xor (X13 and X20 and X32) xor (X13 and X20 and X33) xor (X13 and X22 and X30) xor (X13 and X22 and X32) xor (X13 and X23 and X32) xor (X42) xor (X02 and X42) xor (X00 and X43) xor (X02 and X43) xor (X03 and X42) xor (X00 and X10 and X43) xor (X00 and X12 and X40) xor (X00 and X12 and X42) xor (X00 and X12 and X43) xor (X00 and X13 and X40) xor (X00 and X13 and X42) xor (X02 and X10 and X42) xor (X02 and X10 and X43) xor (X02 and X13 and X40) xor (X02 and X13 and X43) xor (X03 and X10 and X40) xor (X03 and X10 and X42) xor (X03 and X10 and X43) xor (X03 and X12 and X40) xor (X03 and X12 and X42) xor (X03 and X13 and X42) xor (X22 and X42) xor (X20 and X43) xor (X22 and X43) xor (X23 and X42) xor (X00 and X20 and X43) xor (X00 and X22 and X40) xor (X00 and X22 and X42) xor (X00 and X22 and X43) xor (X00 and X23 and X40) xor (X00 and X23 and X42) xor (X02 and X20 and X42) xor (X02 and X20 and X43) xor (X02 and X23 and X40) xor (X02 and X23 and X43) xor (X03 and X20 and X40) xor (X03 and X20 and X42) xor (X03 and X20 and X43) xor (X03 and X22 and X40) xor (X03 and X22 and X42) xor (X03 and X23 and X42) xor (X10 and X20 and X43) xor (X10 and X22 and X40) xor (X10 and X22 and X42) xor (X10 and X22 and X43) xor (X10 and X23 and X40) xor (X10 and X23 and X42) xor (X12 and X20 and X42) xor (X12 and X20 and X43) xor (X12 and X23 and X40) xor (X12 and X23 and X43) xor (X13 and X20 and X40) xor (X13 and X20 and X42) xor (X13 and X20 and X43) xor (X13 and X22 and X40) xor (X13 and X22 and X42) xor (X13 and X23 and X42) xor (X32 and X42) xor (X30 and X43) xor (X32 and X43) xor (X33 and X42) xor (X00 and X30 and X43) xor (X00 and X32 and X40) xor (X00 and X32 and X42) xor (X00 and X32 and X43) xor (X00 and X33 and X40) xor (X00 and X33 and X42) xor (X02 and X30 and X42) xor (X02 and X30 and X43) xor (X02 and X33 and X40) xor (X02 and X33 and X43) xor (X03 and X30 and X40) xor (X03 and X30 and X42) xor (X03 and X30 and X43) xor (X03 and X32 and X40) xor (X03 and X32 and X42) xor (X03 and X33 and X42) xor (X02 and X52) xor (X00 and X53) xor (X02 and X53) xor (X03 and X52) xor (X22 and X52) xor (X20 and X53) xor (X22 and X53) xor (X23 and X52) xor (X10 and X20 and X53) xor (X10 and X22 and X50) xor (X10 and X22 and X52) xor (X10 and X22 and X53) xor (X10 and X23 and X50) xor (X10 and X23 and X52) xor (X12 and X20 and X52) xor (X12 and X20 and X53) xor (X12 and X23 and X50) xor (X12 and X23 and X53) xor (X13 and X20 and X50) xor (X13 and X20 and X52) xor (X13 and X20 and X53) xor (X13 and X22 and X50) xor (X13 and X22 and X52) xor (X13 and X23 and X52) xor (X00 and X30 and X53) xor (X00 and X32 and X50) xor (X00 and X32 and X52) xor (X00 and X32 and X53) xor (X00 and X33 and X50) xor (X00 and X33 and X52) xor (X02 and X30 and X52) xor (X02 and X30 and X53) xor (X02 and X33 and X50) xor (X02 and X33 and X53) xor (X03 and X30 and X50) xor (X03 and X30 and X52) xor (X03 and X30 and X53) xor (X03 and X32 and X50) xor (X03 and X32 and X52) xor (X03 and X33 and X52) xor (X42 and X52) xor (X40 and X53) xor (X42 and X53) xor (X43 and X52) xor (X30 and X40 and X53) xor (X30 and X42 and X50) xor (X30 and X42 and X52) xor (X30 and X42 and X53) xor (X30 and X43 and X50) xor (X30 and X43 and X52) xor (X32 and X40 and X52) xor (X32 and X40 and X53) xor (X32 and X43 and X50) xor (X32 and X43 and X53) xor (X33 and X40 and X50) xor (X33 and X40 and X52) xor (X33 and X40 and X53) xor (X33 and X42 and X50) xor (X33 and X42 and X52) xor (X33 and X43 and X52) xor (X62) xor (X02 and X62) xor (X00 and X63) xor (X02 and X63) xor (X03 and X62) xor (X12 and X62) xor (X10 and X63) xor (X12 and X63) xor (X13 and X62) xor (X32 and X62) xor (X30 and X63) xor (X32 and X63) xor (X33 and X62) xor (X42 and X62) xor (X40 and X63) xor (X42 and X63) xor (X43 and X62) xor (X10 and X40 and X63) xor (X10 and X42 and X60) xor (X10 and X42 and X62) xor (X10 and X42 and X63) xor (X10 and X43 and X60) xor (X10 and X43 and X62) xor (X12 and X40 and X62) xor (X12 and X40 and X63) xor (X12 and X43 and X60) xor (X12 and X43 and X63) xor (X13 and X40 and X60) xor (X13 and X40 and X62) xor (X13 and X40 and X63) xor (X13 and X42 and X60) xor (X13 and X42 and X62) xor (X13 and X43 and X62) xor (X30 and X40 and X63) xor (X30 and X42 and X60) xor (X30 and X42 and X62) xor (X30 and X42 and X63) xor (X30 and X43 and X60) xor (X30 and X43 and X62) xor (X32 and X40 and X62) xor (X32 and X40 and X63) xor (X32 and X43 and X60) xor (X32 and X43 and X63) xor (X33 and X40 and X60) xor (X33 and X40 and X62) xor (X33 and X40 and X63) xor (X33 and X42 and X60) xor (X33 and X42 and X62) xor (X33 and X43 and X62) xor (X10 and X50 and X63) xor (X10 and X52 and X60) xor (X10 and X52 and X62) xor (X10 and X52 and X63) xor (X10 and X53 and X60) xor (X10 and X53 and X62) xor (X12 and X50 and X62) xor (X12 and X50 and X63) xor (X12 and X53 and X60) xor (X12 and X53 and X63) xor (X13 and X50 and X60) xor (X13 and X50 and X62) xor (X13 and X50 and X63) xor (X13 and X52 and X60) xor (X13 and X52 and X62) xor (X13 and X53 and X62) xor (X20 and X50 and X63) xor (X20 and X52 and X60) xor (X20 and X52 and X62) xor (X20 and X52 and X63) xor (X20 and X53 and X60) xor (X20 and X53 and X62) xor (X22 and X50 and X62) xor (X22 and X50 and X63) xor (X22 and X53 and X60) xor (X22 and X53 and X63) xor (X23 and X50 and X60) xor (X23 and X50 and X62) xor (X23 and X50 and X63) xor (X23 and X52 and X60) xor (X23 and X52 and X62) xor (X23 and X53 and X62) xor (X30 and X50 and X63) xor (X30 and X52 and X60) xor (X30 and X52 and X62) xor (X30 and X52 and X63) xor (X30 and X53 and X60) xor (X30 and X53 and X62) xor (X32 and X50 and X62) xor (X32 and X50 and X63) xor (X32 and X53 and X60) xor (X32 and X53 and X63) xor (X33 and X50 and X60) xor (X33 and X50 and X62) xor (X33 and X50 and X63) xor (X33 and X52 and X60) xor (X33 and X52 and X62) xor (X33 and X53 and X62) xor (X00 and X10 and X73) xor (X00 and X12 and X70) xor (X00 and X12 and X72) xor (X00 and X12 and X73) xor (X00 and X13 and X70) xor (X00 and X13 and X72) xor (X02 and X10 and X72) xor (X02 and X10 and X73) xor (X02 and X13 and X70) xor (X02 and X13 and X73) xor (X03 and X10 and X70) xor (X03 and X10 and X72) xor (X03 and X10 and X73) xor (X03 and X12 and X70) xor (X03 and X12 and X72) xor (X03 and X13 and X72) xor (X00 and X20 and X73) xor (X00 and X22 and X70) xor (X00 and X22 and X72) xor (X00 and X22 and X73) xor (X00 and X23 and X70) xor (X00 and X23 and X72) xor (X02 and X20 and X72) xor (X02 and X20 and X73) xor (X02 and X23 and X70) xor (X02 and X23 and X73) xor (X03 and X20 and X70) xor (X03 and X20 and X72) xor (X03 and X20 and X73) xor (X03 and X22 and X70) xor (X03 and X22 and X72) xor (X03 and X23 and X72) xor (X10 and X20 and X73) xor (X10 and X22 and X70) xor (X10 and X22 and X72) xor (X10 and X22 and X73) xor (X10 and X23 and X70) xor (X10 and X23 and X72) xor (X12 and X20 and X72) xor (X12 and X20 and X73) xor (X12 and X23 and X70) xor (X12 and X23 and X73) xor (X13 and X20 and X70) xor (X13 and X20 and X72) xor (X13 and X20 and X73) xor (X13 and X22 and X70) xor (X13 and X22 and X72) xor (X13 and X23 and X72) xor (X32 and X72) xor (X30 and X73) xor (X32 and X73) xor (X33 and X72) xor (X10 and X30 and X73) xor (X10 and X32 and X70) xor (X10 and X32 and X72) xor (X10 and X32 and X73) xor (X10 and X33 and X70) xor (X10 and X33 and X72) xor (X12 and X30 and X72) xor (X12 and X30 and X73) xor (X12 and X33 and X70) xor (X12 and X33 and X73) xor (X13 and X30 and X70) xor (X13 and X30 and X72) xor (X13 and X30 and X73) xor (X13 and X32 and X70) xor (X13 and X32 and X72) xor (X13 and X33 and X72) xor (X42 and X72) xor (X40 and X73) xor (X42 and X73) xor (X43 and X72) xor (X00 and X40 and X73) xor (X00 and X42 and X70) xor (X00 and X42 and X72) xor (X00 and X42 and X73) xor (X00 and X43 and X70) xor (X00 and X43 and X72) xor (X02 and X40 and X72) xor (X02 and X40 and X73) xor (X02 and X43 and X70) xor (X02 and X43 and X73) xor (X03 and X40 and X70) xor (X03 and X40 and X72) xor (X03 and X40 and X73) xor (X03 and X42 and X70) xor (X03 and X42 and X72) xor (X03 and X43 and X72) xor (X10 and X40 and X73) xor (X10 and X42 and X70) xor (X10 and X42 and X72) xor (X10 and X42 and X73) xor (X10 and X43 and X70) xor (X10 and X43 and X72) xor (X12 and X40 and X72) xor (X12 and X40 and X73) xor (X12 and X43 and X70) xor (X12 and X43 and X73) xor (X13 and X40 and X70) xor (X13 and X40 and X72) xor (X13 and X40 and X73) xor (X13 and X42 and X70) xor (X13 and X42 and X72) xor (X13 and X43 and X72) xor (X20 and X40 and X73) xor (X20 and X42 and X70) xor (X20 and X42 and X72) xor (X20 and X42 and X73) xor (X20 and X43 and X70) xor (X20 and X43 and X72) xor (X22 and X40 and X72) xor (X22 and X40 and X73) xor (X22 and X43 and X70) xor (X22 and X43 and X73) xor (X23 and X40 and X70) xor (X23 and X40 and X72) xor (X23 and X40 and X73) xor (X23 and X42 and X70) xor (X23 and X42 and X72) xor (X23 and X43 and X72) xor (X52 and X72) xor (X50 and X73) xor (X52 and X73) xor (X53 and X72) xor (X00 and X50 and X73) xor (X00 and X52 and X70) xor (X00 and X52 and X72) xor (X00 and X52 and X73) xor (X00 and X53 and X70) xor (X00 and X53 and X72) xor (X02 and X50 and X72) xor (X02 and X50 and X73) xor (X02 and X53 and X70) xor (X02 and X53 and X73) xor (X03 and X50 and X70) xor (X03 and X50 and X72) xor (X03 and X50 and X73) xor (X03 and X52 and X70) xor (X03 and X52 and X72) xor (X03 and X53 and X72) xor (X62 and X72) xor (X60 and X73) xor (X62 and X73) xor (X63 and X72) xor (X00 and X60 and X73) xor (X00 and X62 and X70) xor (X00 and X62 and X72) xor (X00 and X62 and X73) xor (X00 and X63 and X70) xor (X00 and X63 and X72) xor (X02 and X60 and X72) xor (X02 and X60 and X73) xor (X02 and X63 and X70) xor (X02 and X63 and X73) xor (X03 and X60 and X70) xor (X03 and X60 and X72) xor (X03 and X60 and X73) xor (X03 and X62 and X70) xor (X03 and X62 and X72) xor (X03 and X63 and X72) xor (X30 and X60 and X73) xor (X30 and X62 and X70) xor (X30 and X62 and X72) xor (X30 and X62 and X73) xor (X30 and X63 and X70) xor (X30 and X63 and X72) xor (X32 and X60 and X72) xor (X32 and X60 and X73) xor (X32 and X63 and X70) xor (X32 and X63 and X73) xor (X33 and X60 and X70) xor (X33 and X60 and X72) xor (X33 and X60 and X73) xor (X33 and X62 and X70) xor (X33 and X62 and X72) xor (X33 and X63 and X72));
    F63  <= ((X13) xor (X23) xor (X13 and X23) xor (X13 and X20) xor (X13 and X21) xor (X11 and X20) xor (X00 and X10 and X21) xor (X00 and X11 and X20) xor (X00 and X11 and X23) xor (X00 and X13 and X21) xor (X00 and X13 and X23) xor (X0_1 and X10 and X21) xor (X0_1 and X10 and X23) xor (X0_1 and X11 and X23) xor (X0_1 and X13 and X20) xor (X0_1 and X13 and X21) xor (X0_1 and X13 and X23) xor (X03 and X10 and X21) xor (X03 and X11 and X20) xor (X03 and X11 and X21) xor (X03 and X11 and X23) xor (X03 and X13 and X20) xor (X03 and X33) xor (X03 and X30) xor (X03 and X31) xor (X0_1 and X30) xor (X23 and X33) xor (X23 and X30) xor (X23 and X31) xor (X21 and X30) xor (X00 and X20 and X31) xor (X00 and X21 and X30) xor (X00 and X21 and X33) xor (X00 and X23 and X31) xor (X00 and X23 and X33) xor (X0_1 and X20 and X31) xor (X0_1 and X20 and X33) xor (X0_1 and X21 and X33) xor (X0_1 and X23 and X30) xor (X0_1 and X23 and X31) xor (X0_1 and X23 and X33) xor (X03 and X20 and X31) xor (X03 and X21 and X30) xor (X03 and X21 and X31) xor (X03 and X21 and X33) xor (X03 and X23 and X30) xor (X10 and X20 and X31) xor (X10 and X21 and X30) xor (X10 and X21 and X33) xor (X10 and X23 and X31) xor (X10 and X23 and X33) xor (X11 and X20 and X31) xor (X11 and X20 and X33) xor (X11 and X21 and X33) xor (X11 and X23 and X30) xor (X11 and X23 and X31) xor (X11 and X23 and X33) xor (X13 and X20 and X31) xor (X13 and X21 and X30) xor (X13 and X21 and X31) xor (X13 and X21 and X33) xor (X13 and X23 and X30) xor (X43) xor (X03 and X43) xor (X03 and X40) xor (X03 and X41) xor (X0_1 and X40) xor (X00 and X10 and X41) xor (X00 and X11 and X40) xor (X00 and X11 and X43) xor (X00 and X13 and X41) xor (X00 and X13 and X43) xor (X0_1 and X10 and X41) xor (X0_1 and X10 and X43) xor (X0_1 and X11 and X43) xor (X0_1 and X13 and X40) xor (X0_1 and X13 and X41) xor (X0_1 and X13 and X43) xor (X03 and X10 and X41) xor (X03 and X11 and X40) xor (X03 and X11 and X41) xor (X03 and X11 and X43) xor (X03 and X13 and X40) xor (X23 and X43) xor (X23 and X40) xor (X23 and X41) xor (X21 and X40) xor (X00 and X20 and X41) xor (X00 and X21 and X40) xor (X00 and X21 and X43) xor (X00 and X23 and X41) xor (X00 and X23 and X43) xor (X0_1 and X20 and X41) xor (X0_1 and X20 and X43) xor (X0_1 and X21 and X43) xor (X0_1 and X23 and X40) xor (X0_1 and X23 and X41) xor (X0_1 and X23 and X43) xor (X03 and X20 and X41) xor (X03 and X21 and X40) xor (X03 and X21 and X41) xor (X03 and X21 and X43) xor (X03 and X23 and X40) xor (X10 and X20 and X41) xor (X10 and X21 and X40) xor (X10 and X21 and X43) xor (X10 and X23 and X41) xor (X10 and X23 and X43) xor (X11 and X20 and X41) xor (X11 and X20 and X43) xor (X11 and X21 and X43) xor (X11 and X23 and X40) xor (X11 and X23 and X41) xor (X11 and X23 and X43) xor (X13 and X20 and X41) xor (X13 and X21 and X40) xor (X13 and X21 and X41) xor (X13 and X21 and X43) xor (X13 and X23 and X40) xor (X33 and X43) xor (X33 and X40) xor (X33 and X41) xor (X31 and X40) xor (X00 and X30 and X41) xor (X00 and X31 and X40) xor (X00 and X31 and X43) xor (X00 and X33 and X41) xor (X00 and X33 and X43) xor (X0_1 and X30 and X41) xor (X0_1 and X30 and X43) xor (X0_1 and X31 and X43) xor (X0_1 and X33 and X40) xor (X0_1 and X33 and X41) xor (X0_1 and X33 and X43) xor (X03 and X30 and X41) xor (X03 and X31 and X40) xor (X03 and X31 and X41) xor (X03 and X31 and X43) xor (X03 and X33 and X40) xor (X03 and X53) xor (X03 and X50) xor (X03 and X51) xor (X0_1 and X50) xor (X23 and X53) xor (X23 and X50) xor (X23 and X51) xor (X21 and X50) xor (X10 and X20 and X51) xor (X10 and X21 and X50) xor (X10 and X21 and X53) xor (X10 and X23 and X51) xor (X10 and X23 and X53) xor (X11 and X20 and X51) xor (X11 and X20 and X53) xor (X11 and X21 and X53) xor (X11 and X23 and X50) xor (X11 and X23 and X51) xor (X11 and X23 and X53) xor (X13 and X20 and X51) xor (X13 and X21 and X50) xor (X13 and X21 and X51) xor (X13 and X21 and X53) xor (X13 and X23 and X50) xor (X00 and X30 and X51) xor (X00 and X31 and X50) xor (X00 and X31 and X53) xor (X00 and X33 and X51) xor (X00 and X33 and X53) xor (X0_1 and X30 and X51) xor (X0_1 and X30 and X53) xor (X0_1 and X31 and X53) xor (X0_1 and X33 and X50) xor (X0_1 and X33 and X51) xor (X0_1 and X33 and X53) xor (X03 and X30 and X51) xor (X03 and X31 and X50) xor (X03 and X31 and X51) xor (X03 and X31 and X53) xor (X03 and X33 and X50) xor (X43 and X53) xor (X43 and X50) xor (X43 and X51) xor (X41 and X50) xor (X30 and X40 and X51) xor (X30 and X41 and X50) xor (X30 and X41 and X53) xor (X30 and X43 and X51) xor (X30 and X43 and X53) xor (X31 and X40 and X51) xor (X31 and X40 and X53) xor (X31 and X41 and X53) xor (X31 and X43 and X50) xor (X31 and X43 and X51) xor (X31 and X43 and X53) xor (X33 and X40 and X51) xor (X33 and X41 and X50) xor (X33 and X41 and X51) xor (X33 and X41 and X53) xor (X33 and X43 and X50) xor (X63) xor (X03 and X63) xor (X03 and X60) xor (X03 and X61) xor (X0_1 and X60) xor (X13 and X63) xor (X13 and X60) xor (X13 and X61) xor (X11 and X60) xor (X33 and X63) xor (X33 and X60) xor (X33 and X61) xor (X31 and X60) xor (X43 and X63) xor (X43 and X60) xor (X43 and X61) xor (X41 and X60) xor (X10 and X40 and X61) xor (X10 and X41 and X60) xor (X10 and X41 and X63) xor (X10 and X43 and X61) xor (X10 and X43 and X63) xor (X11 and X40 and X61) xor (X11 and X40 and X63) xor (X11 and X41 and X63) xor (X11 and X43 and X60) xor (X11 and X43 and X61) xor (X11 and X43 and X63) xor (X13 and X40 and X61) xor (X13 and X41 and X60) xor (X13 and X41 and X61) xor (X13 and X41 and X63) xor (X13 and X43 and X60) xor (X30 and X40 and X61) xor (X30 and X41 and X60) xor (X30 and X41 and X63) xor (X30 and X43 and X61) xor (X30 and X43 and X63) xor (X31 and X40 and X61) xor (X31 and X40 and X63) xor (X31 and X41 and X63) xor (X31 and X43 and X60) xor (X31 and X43 and X61) xor (X31 and X43 and X63) xor (X33 and X40 and X61) xor (X33 and X41 and X60) xor (X33 and X41 and X61) xor (X33 and X41 and X63) xor (X33 and X43 and X60) xor (X10 and X50 and X61) xor (X10 and X51 and X60) xor (X10 and X51 and X63) xor (X10 and X53 and X61) xor (X10 and X53 and X63) xor (X11 and X50 and X61) xor (X11 and X50 and X63) xor (X11 and X51 and X63) xor (X11 and X53 and X60) xor (X11 and X53 and X61) xor (X11 and X53 and X63) xor (X13 and X50 and X61) xor (X13 and X51 and X60) xor (X13 and X51 and X61) xor (X13 and X51 and X63) xor (X13 and X53 and X60) xor (X20 and X50 and X61) xor (X20 and X51 and X60) xor (X20 and X51 and X63) xor (X20 and X53 and X61) xor (X20 and X53 and X63) xor (X21 and X50 and X61) xor (X21 and X50 and X63) xor (X21 and X51 and X63) xor (X21 and X53 and X60) xor (X21 and X53 and X61) xor (X21 and X53 and X63) xor (X23 and X50 and X61) xor (X23 and X51 and X60) xor (X23 and X51 and X61) xor (X23 and X51 and X63) xor (X23 and X53 and X60) xor (X30 and X50 and X61) xor (X30 and X51 and X60) xor (X30 and X51 and X63) xor (X30 and X53 and X61) xor (X30 and X53 and X63) xor (X31 and X50 and X61) xor (X31 and X50 and X63) xor (X31 and X51 and X63) xor (X31 and X53 and X60) xor (X31 and X53 and X61) xor (X31 and X53 and X63) xor (X33 and X50 and X61) xor (X33 and X51 and X60) xor (X33 and X51 and X61) xor (X33 and X51 and X63) xor (X33 and X53 and X60) xor (X00 and X10 and X71) xor (X00 and X11 and X70) xor (X00 and X11 and X73) xor (X00 and X13 and X71) xor (X00 and X13 and X73) xor (X0_1 and X10 and X71) xor (X0_1 and X10 and X73) xor (X0_1 and X11 and X73) xor (X0_1 and X13 and X70) xor (X0_1 and X13 and X71) xor (X0_1 and X13 and X73) xor (X03 and X10 and X71) xor (X03 and X11 and X70) xor (X03 and X11 and X71) xor (X03 and X11 and X73) xor (X03 and X13 and X70) xor (X00 and X20 and X71) xor (X00 and X21 and X70) xor (X00 and X21 and X73) xor (X00 and X23 and X71) xor (X00 and X23 and X73) xor (X0_1 and X20 and X71) xor (X0_1 and X20 and X73) xor (X0_1 and X21 and X73) xor (X0_1 and X23 and X70) xor (X0_1 and X23 and X71) xor (X0_1 and X23 and X73) xor (X03 and X20 and X71) xor (X03 and X21 and X70) xor (X03 and X21 and X71) xor (X03 and X21 and X73) xor (X03 and X23 and X70) xor (X10 and X20 and X71) xor (X10 and X21 and X70) xor (X10 and X21 and X73) xor (X10 and X23 and X71) xor (X10 and X23 and X73) xor (X11 and X20 and X71) xor (X11 and X20 and X73) xor (X11 and X21 and X73) xor (X11 and X23 and X70) xor (X11 and X23 and X71) xor (X11 and X23 and X73) xor (X13 and X20 and X71) xor (X13 and X21 and X70) xor (X13 and X21 and X71) xor (X13 and X21 and X73) xor (X13 and X23 and X70) xor (X33 and X73) xor (X33 and X70) xor (X33 and X71) xor (X31 and X70) xor (X10 and X30 and X71) xor (X10 and X31 and X70) xor (X10 and X31 and X73) xor (X10 and X33 and X71) xor (X10 and X33 and X73) xor (X11 and X30 and X71) xor (X11 and X30 and X73) xor (X11 and X31 and X73) xor (X11 and X33 and X70) xor (X11 and X33 and X71) xor (X11 and X33 and X73) xor (X13 and X30 and X71) xor (X13 and X31 and X70) xor (X13 and X31 and X71) xor (X13 and X31 and X73) xor (X13 and X33 and X70) xor (X43 and X73) xor (X43 and X70) xor (X43 and X71) xor (X41 and X70) xor (X00 and X40 and X71) xor (X00 and X41 and X70) xor (X00 and X41 and X73) xor (X00 and X43 and X71) xor (X00 and X43 and X73) xor (X0_1 and X40 and X71) xor (X0_1 and X40 and X73) xor (X0_1 and X41 and X73) xor (X0_1 and X43 and X70) xor (X0_1 and X43 and X71) xor (X0_1 and X43 and X73) xor (X03 and X40 and X71) xor (X03 and X41 and X70) xor (X03 and X41 and X71) xor (X03 and X41 and X73) xor (X03 and X43 and X70) xor (X10 and X40 and X71) xor (X10 and X41 and X70) xor (X10 and X41 and X73) xor (X10 and X43 and X71) xor (X10 and X43 and X73) xor (X11 and X40 and X71) xor (X11 and X40 and X73) xor (X11 and X41 and X73) xor (X11 and X43 and X70) xor (X11 and X43 and X71) xor (X11 and X43 and X73) xor (X13 and X40 and X71) xor (X13 and X41 and X70) xor (X13 and X41 and X71) xor (X13 and X41 and X73) xor (X13 and X43 and X70) xor (X20 and X40 and X71) xor (X20 and X41 and X70) xor (X20 and X41 and X73) xor (X20 and X43 and X71) xor (X20 and X43 and X73) xor (X21 and X40 and X71) xor (X21 and X40 and X73) xor (X21 and X41 and X73) xor (X21 and X43 and X70) xor (X21 and X43 and X71) xor (X21 and X43 and X73) xor (X23 and X40 and X71) xor (X23 and X41 and X70) xor (X23 and X41 and X71) xor (X23 and X41 and X73) xor (X23 and X43 and X70) xor (X53 and X73) xor (X53 and X70) xor (X53 and X71) xor (X51 and X70) xor (X00 and X50 and X71) xor (X00 and X51 and X70) xor (X00 and X51 and X73) xor (X00 and X53 and X71) xor (X00 and X53 and X73) xor (X0_1 and X50 and X71) xor (X0_1 and X50 and X73) xor (X0_1 and X51 and X73) xor (X0_1 and X53 and X70) xor (X0_1 and X53 and X71) xor (X0_1 and X53 and X73) xor (X03 and X50 and X71) xor (X03 and X51 and X70) xor (X03 and X51 and X71) xor (X03 and X51 and X73) xor (X03 and X53 and X70) xor (X63 and X73) xor (X63 and X70) xor (X63 and X71) xor (X61 and X70) xor (X00 and X60 and X71) xor (X00 and X61 and X70) xor (X00 and X61 and X73) xor (X00 and X63 and X71) xor (X00 and X63 and X73) xor (X0_1 and X60 and X71) xor (X0_1 and X60 and X73) xor (X0_1 and X61 and X73) xor (X0_1 and X63 and X70) xor (X0_1 and X63 and X71) xor (X0_1 and X63 and X73) xor (X03 and X60 and X71) xor (X03 and X61 and X70) xor (X03 and X61 and X71) xor (X03 and X61 and X73) xor (X03 and X63 and X70) xor (X30 and X60 and X71) xor (X30 and X61 and X70) xor (X30 and X61 and X73) xor (X30 and X63 and X71) xor (X30 and X63 and X73) xor (X31 and X60 and X71) xor (X31 and X60 and X73) xor (X31 and X61 and X73) xor (X31 and X63 and X70) xor (X31 and X63 and X71) xor (X31 and X63 and X73) xor (X33 and X60 and X71) xor (X33 and X61 and X70) xor (X33 and X61 and X71) xor (X33 and X61 and X73) xor (X33 and X63 and X70));
    F70  <= ((X10) xor (X10 and X30) xor (X10 and X31) xor (X12 and X30) xor (X10 and X32) xor (X00 and X10 and X30) xor (X00 and X10 and X32) xor (X00 and X11 and X31) xor (X00 and X11 and X32) xor (X00 and X12 and X31) xor (X0_1 and X10 and X30) xor (X0_1 and X10 and X32) xor (X0_1 and X11 and X30) xor (X0_1 and X12 and X30) xor (X0_1 and X12 and X31) xor (X02 and X10 and X30) xor (X02 and X10 and X31) xor (X02 and X11 and X30) xor (X02 and X11 and X31) xor (X02 and X12 and X30) xor (X02 and X12 and X32) xor (X20 and X30) xor (X20 and X31) xor (X22 and X30) xor (X20 and X32) xor (X40) xor (X10 and X40) xor (X10 and X41) xor (X12 and X40) xor (X10 and X42) xor (X20 and X40) xor (X20 and X41) xor (X22 and X40) xor (X20 and X42) xor (X00 and X20 and X40) xor (X00 and X20 and X42) xor (X00 and X21 and X41) xor (X00 and X21 and X42) xor (X00 and X22 and X41) xor (X0_1 and X20 and X40) xor (X0_1 and X20 and X42) xor (X0_1 and X21 and X40) xor (X0_1 and X22 and X40) xor (X0_1 and X22 and X41) xor (X02 and X20 and X40) xor (X02 and X20 and X41) xor (X02 and X21 and X40) xor (X02 and X21 and X41) xor (X02 and X22 and X40) xor (X02 and X22 and X42) xor (X30 and X40) xor (X30 and X41) xor (X32 and X40) xor (X30 and X42) xor (X00 and X50) xor (X00 and X51) xor (X02 and X50) xor (X00 and X52) xor (X20 and X50) xor (X20 and X51) xor (X22 and X50) xor (X20 and X52) xor (X00 and X20 and X50) xor (X00 and X20 and X52) xor (X00 and X21 and X51) xor (X00 and X21 and X52) xor (X00 and X22 and X51) xor (X0_1 and X20 and X50) xor (X0_1 and X20 and X52) xor (X0_1 and X21 and X50) xor (X0_1 and X22 and X50) xor (X0_1 and X22 and X51) xor (X02 and X20 and X50) xor (X02 and X20 and X51) xor (X02 and X21 and X50) xor (X02 and X21 and X51) xor (X02 and X22 and X50) xor (X02 and X22 and X52) xor (X30 and X50) xor (X30 and X51) xor (X32 and X50) xor (X30 and X52) xor (X00 and X30 and X50) xor (X00 and X30 and X52) xor (X00 and X31 and X51) xor (X00 and X31 and X52) xor (X00 and X32 and X51) xor (X0_1 and X30 and X50) xor (X0_1 and X30 and X52) xor (X0_1 and X31 and X50) xor (X0_1 and X32 and X50) xor (X0_1 and X32 and X51) xor (X02 and X30 and X50) xor (X02 and X30 and X51) xor (X02 and X31 and X50) xor (X02 and X31 and X51) xor (X02 and X32 and X50) xor (X02 and X32 and X52) xor (X10 and X30 and X50) xor (X10 and X30 and X52) xor (X10 and X31 and X51) xor (X10 and X31 and X52) xor (X10 and X32 and X51) xor (X11 and X30 and X50) xor (X11 and X30 and X52) xor (X11 and X31 and X50) xor (X11 and X32 and X50) xor (X11 and X32 and X51) xor (X12 and X30 and X50) xor (X12 and X30 and X51) xor (X12 and X31 and X50) xor (X12 and X31 and X51) xor (X12 and X32 and X50) xor (X12 and X32 and X52) xor (X40 and X50) xor (X40 and X51) xor (X42 and X50) xor (X40 and X52) xor (X00 and X40 and X50) xor (X00 and X40 and X52) xor (X00 and X41 and X51) xor (X00 and X41 and X52) xor (X00 and X42 and X51) xor (X0_1 and X40 and X50) xor (X0_1 and X40 and X52) xor (X0_1 and X41 and X50) xor (X0_1 and X42 and X50) xor (X0_1 and X42 and X51) xor (X02 and X40 and X50) xor (X02 and X40 and X51) xor (X02 and X41 and X50) xor (X02 and X41 and X51) xor (X02 and X42 and X50) xor (X02 and X42 and X52) xor (X10 and X40 and X50) xor (X10 and X40 and X52) xor (X10 and X41 and X51) xor (X10 and X41 and X52) xor (X10 and X42 and X51) xor (X11 and X40 and X50) xor (X11 and X40 and X52) xor (X11 and X41 and X50) xor (X11 and X42 and X50) xor (X11 and X42 and X51) xor (X12 and X40 and X50) xor (X12 and X40 and X51) xor (X12 and X41 and X50) xor (X12 and X41 and X51) xor (X12 and X42 and X50) xor (X12 and X42 and X52) xor (X30 and X40 and X50) xor (X30 and X40 and X52) xor (X30 and X41 and X51) xor (X30 and X41 and X52) xor (X30 and X42 and X51) xor (X31 and X40 and X50) xor (X31 and X40 and X52) xor (X31 and X41 and X50) xor (X31 and X42 and X50) xor (X31 and X42 and X51) xor (X32 and X40 and X50) xor (X32 and X40 and X51) xor (X32 and X41 and X50) xor (X32 and X41 and X51) xor (X32 and X42 and X50) xor (X32 and X42 and X52) xor (X00 and X60) xor (X00 and X61) xor (X02 and X60) xor (X00 and X62) xor (X10 and X60) xor (X10 and X61) xor (X12 and X60) xor (X10 and X62) xor (X20 and X60) xor (X20 and X61) xor (X22 and X60) xor (X20 and X62) xor (X00 and X20 and X60) xor (X00 and X20 and X62) xor (X00 and X21 and X61) xor (X00 and X21 and X62) xor (X00 and X22 and X61) xor (X0_1 and X20 and X60) xor (X0_1 and X20 and X62) xor (X0_1 and X21 and X60) xor (X0_1 and X22 and X60) xor (X0_1 and X22 and X61) xor (X02 and X20 and X60) xor (X02 and X20 and X61) xor (X02 and X21 and X60) xor (X02 and X21 and X61) xor (X02 and X22 and X60) xor (X02 and X22 and X62) xor (X00 and X40 and X60) xor (X00 and X40 and X62) xor (X00 and X41 and X61) xor (X00 and X41 and X62) xor (X00 and X42 and X61) xor (X0_1 and X40 and X60) xor (X0_1 and X40 and X62) xor (X0_1 and X41 and X60) xor (X0_1 and X42 and X60) xor (X0_1 and X42 and X61) xor (X02 and X40 and X60) xor (X02 and X40 and X61) xor (X02 and X41 and X60) xor (X02 and X41 and X61) xor (X02 and X42 and X60) xor (X02 and X42 and X62) xor (X10 and X40 and X60) xor (X10 and X40 and X62) xor (X10 and X41 and X61) xor (X10 and X41 and X62) xor (X10 and X42 and X61) xor (X11 and X40 and X60) xor (X11 and X40 and X62) xor (X11 and X41 and X60) xor (X11 and X42 and X60) xor (X11 and X42 and X61) xor (X12 and X40 and X60) xor (X12 and X40 and X61) xor (X12 and X41 and X60) xor (X12 and X41 and X61) xor (X12 and X42 and X60) xor (X12 and X42 and X62) xor (X20 and X40 and X60) xor (X20 and X40 and X62) xor (X20 and X41 and X61) xor (X20 and X41 and X62) xor (X20 and X42 and X61) xor (X21 and X40 and X60) xor (X21 and X40 and X62) xor (X21 and X41 and X60) xor (X21 and X42 and X60) xor (X21 and X42 and X61) xor (X22 and X40 and X60) xor (X22 and X40 and X61) xor (X22 and X41 and X60) xor (X22 and X41 and X61) xor (X22 and X42 and X60) xor (X22 and X42 and X62) xor (X00 and X50 and X60) xor (X00 and X50 and X62) xor (X00 and X51 and X61) xor (X00 and X51 and X62) xor (X00 and X52 and X61) xor (X0_1 and X50 and X60) xor (X0_1 and X50 and X62) xor (X0_1 and X51 and X60) xor (X0_1 and X52 and X60) xor (X0_1 and X52 and X61) xor (X02 and X50 and X60) xor (X02 and X50 and X61) xor (X02 and X51 and X60) xor (X02 and X51 and X61) xor (X02 and X52 and X60) xor (X02 and X52 and X62) xor (X10 and X50 and X60) xor (X10 and X50 and X62) xor (X10 and X51 and X61) xor (X10 and X51 and X62) xor (X10 and X52 and X61) xor (X11 and X50 and X60) xor (X11 and X50 and X62) xor (X11 and X51 and X60) xor (X11 and X52 and X60) xor (X11 and X52 and X61) xor (X12 and X50 and X60) xor (X12 and X50 and X61) xor (X12 and X51 and X60) xor (X12 and X51 and X61) xor (X12 and X52 and X60) xor (X12 and X52 and X62) xor (X20 and X50 and X60) xor (X20 and X50 and X62) xor (X20 and X51 and X61) xor (X20 and X51 and X62) xor (X20 and X52 and X61) xor (X21 and X50 and X60) xor (X21 and X50 and X62) xor (X21 and X51 and X60) xor (X21 and X52 and X60) xor (X21 and X52 and X61) xor (X22 and X50 and X60) xor (X22 and X50 and X61) xor (X22 and X51 and X60) xor (X22 and X51 and X61) xor (X22 and X52 and X60) xor (X22 and X52 and X62) xor (X30 and X50 and X60) xor (X30 and X50 and X62) xor (X30 and X51 and X61) xor (X30 and X51 and X62) xor (X30 and X52 and X61) xor (X31 and X50 and X60) xor (X31 and X50 and X62) xor (X31 and X51 and X60) xor (X31 and X52 and X60) xor (X31 and X52 and X61) xor (X32 and X50 and X60) xor (X32 and X50 and X61) xor (X32 and X51 and X60) xor (X32 and X51 and X61) xor (X32 and X52 and X60) xor (X32 and X52 and X62) xor (X40 and X50 and X60) xor (X40 and X50 and X62) xor (X40 and X51 and X61) xor (X40 and X51 and X62) xor (X40 and X52 and X61) xor (X41 and X50 and X60) xor (X41 and X50 and X62) xor (X41 and X51 and X60) xor (X41 and X52 and X60) xor (X41 and X52 and X61) xor (X42 and X50 and X60) xor (X42 and X50 and X61) xor (X42 and X51 and X60) xor (X42 and X51 and X61) xor (X42 and X52 and X60) xor (X42 and X52 and X62) xor (X70) xor (X00 and X10 and X70) xor (X00 and X10 and X72) xor (X00 and X11 and X71) xor (X00 and X11 and X72) xor (X00 and X12 and X71) xor (X0_1 and X10 and X70) xor (X0_1 and X10 and X72) xor (X0_1 and X11 and X70) xor (X0_1 and X12 and X70) xor (X0_1 and X12 and X71) xor (X02 and X10 and X70) xor (X02 and X10 and X71) xor (X02 and X11 and X70) xor (X02 and X11 and X71) xor (X02 and X12 and X70) xor (X02 and X12 and X72) xor (X20 and X70) xor (X20 and X71) xor (X22 and X70) xor (X20 and X72) xor (X00 and X20 and X70) xor (X00 and X20 and X72) xor (X00 and X21 and X71) xor (X00 and X21 and X72) xor (X00 and X22 and X71) xor (X0_1 and X20 and X70) xor (X0_1 and X20 and X72) xor (X0_1 and X21 and X70) xor (X0_1 and X22 and X70) xor (X0_1 and X22 and X71) xor (X02 and X20 and X70) xor (X02 and X20 and X71) xor (X02 and X21 and X70) xor (X02 and X21 and X71) xor (X02 and X22 and X70) xor (X02 and X22 and X72) xor (X40 and X70) xor (X40 and X71) xor (X42 and X70) xor (X40 and X72) xor (X20 and X40 and X70) xor (X20 and X40 and X72) xor (X20 and X41 and X71) xor (X20 and X41 and X72) xor (X20 and X42 and X71) xor (X21 and X40 and X70) xor (X21 and X40 and X72) xor (X21 and X41 and X70) xor (X21 and X42 and X70) xor (X21 and X42 and X71) xor (X22 and X40 and X70) xor (X22 and X40 and X71) xor (X22 and X41 and X70) xor (X22 and X41 and X71) xor (X22 and X42 and X70) xor (X22 and X42 and X72) xor (X20 and X50 and X70) xor (X20 and X50 and X72) xor (X20 and X51 and X71) xor (X20 and X51 and X72) xor (X20 and X52 and X71) xor (X21 and X50 and X70) xor (X21 and X50 and X72) xor (X21 and X51 and X70) xor (X21 and X52 and X70) xor (X21 and X52 and X71) xor (X22 and X50 and X70) xor (X22 and X50 and X71) xor (X22 and X51 and X70) xor (X22 and X51 and X71) xor (X22 and X52 and X70) xor (X22 and X52 and X72) xor (X60 and X70) xor (X60 and X71) xor (X62 and X70) xor (X60 and X72) xor (X00 and X60 and X70) xor (X00 and X60 and X72) xor (X00 and X61 and X71) xor (X00 and X61 and X72) xor (X00 and X62 and X71) xor (X0_1 and X60 and X70) xor (X0_1 and X60 and X72) xor (X0_1 and X61 and X70) xor (X0_1 and X62 and X70) xor (X0_1 and X62 and X71) xor (X02 and X60 and X70) xor (X02 and X60 and X71) xor (X02 and X61 and X70) xor (X02 and X61 and X71) xor (X02 and X62 and X70) xor (X02 and X62 and X72) xor (X30 and X60 and X70) xor (X30 and X60 and X72) xor (X30 and X61 and X71) xor (X30 and X61 and X72) xor (X30 and X62 and X71) xor (X31 and X60 and X70) xor (X31 and X60 and X72) xor (X31 and X61 and X70) xor (X31 and X62 and X70) xor (X31 and X62 and X71) xor (X32 and X60 and X70) xor (X32 and X60 and X71) xor (X32 and X61 and X70) xor (X32 and X61 and X71) xor (X32 and X62 and X70) xor (X32 and X62 and X72) xor (X40 and X60 and X70) xor (X40 and X60 and X72) xor (X40 and X61 and X71) xor (X40 and X61 and X72) xor (X40 and X62 and X71) xor (X41 and X60 and X70) xor (X41 and X60 and X72) xor (X41 and X61 and X70) xor (X41 and X62 and X70) xor (X41 and X62 and X71) xor (X42 and X60 and X70) xor (X42 and X60 and X71) xor (X42 and X61 and X70) xor (X42 and X61 and X71) xor (X42 and X62 and X70) xor (X42 and X62 and X72) xor (X50 and X60 and X70) xor (X50 and X60 and X72) xor (X50 and X61 and X71) xor (X50 and X61 and X72) xor (X50 and X62 and X71) xor (X51 and X60 and X70) xor (X51 and X60 and X72) xor (X51 and X61 and X70) xor (X51 and X62 and X70) xor (X51 and X62 and X71) xor (X52 and X60 and X70) xor (X52 and X60 and X71) xor (X52 and X61 and X70) xor (X52 and X61 and X71) xor (X52 and X62 and X70) xor (X52 and X62 and X72));
    F71  <= ((X11) xor (X11 and X31) xor (X11 and X32) xor (X12 and X31) xor (X11 and X33) xor (X0_1 and X11 and X31) xor (X0_1 and X11 and X32) xor (X0_1 and X12 and X32) xor (X0_1 and X12 and X33) xor (X0_1 and X13 and X32) xor (X02 and X11 and X32) xor (X02 and X11 and X33) xor (X02 and X12 and X31) xor (X02 and X12 and X33) xor (X02 and X13 and X31) xor (X02 and X13 and X32) xor (X03 and X11 and X32) xor (X03 and X12 and X31) xor (X03 and X12 and X33) xor (X03 and X13 and X31) xor (X03 and X13 and X33) xor (X21 and X31) xor (X21 and X32) xor (X22 and X31) xor (X21 and X33) xor (X41) xor (X11 and X41) xor (X11 and X42) xor (X12 and X41) xor (X11 and X43) xor (X21 and X41) xor (X21 and X42) xor (X22 and X41) xor (X21 and X43) xor (X0_1 and X21 and X41) xor (X0_1 and X21 and X42) xor (X0_1 and X22 and X42) xor (X0_1 and X22 and X43) xor (X0_1 and X23 and X42) xor (X02 and X21 and X42) xor (X02 and X21 and X43) xor (X02 and X22 and X41) xor (X02 and X22 and X43) xor (X02 and X23 and X41) xor (X02 and X23 and X42) xor (X03 and X21 and X42) xor (X03 and X22 and X41) xor (X03 and X22 and X43) xor (X03 and X23 and X41) xor (X03 and X23 and X43) xor (X31 and X41) xor (X31 and X42) xor (X32 and X41) xor (X31 and X43) xor (X0_1 and X51) xor (X0_1 and X52) xor (X02 and X51) xor (X0_1 and X53) xor (X21 and X51) xor (X21 and X52) xor (X22 and X51) xor (X21 and X53) xor (X0_1 and X21 and X51) xor (X0_1 and X21 and X52) xor (X0_1 and X22 and X52) xor (X0_1 and X22 and X53) xor (X0_1 and X23 and X52) xor (X02 and X21 and X52) xor (X02 and X21 and X53) xor (X02 and X22 and X51) xor (X02 and X22 and X53) xor (X02 and X23 and X51) xor (X02 and X23 and X52) xor (X03 and X21 and X52) xor (X03 and X22 and X51) xor (X03 and X22 and X53) xor (X03 and X23 and X51) xor (X03 and X23 and X53) xor (X31 and X51) xor (X31 and X52) xor (X32 and X51) xor (X31 and X53) xor (X0_1 and X31 and X51) xor (X0_1 and X31 and X52) xor (X0_1 and X32 and X52) xor (X0_1 and X32 and X53) xor (X0_1 and X33 and X52) xor (X02 and X31 and X52) xor (X02 and X31 and X53) xor (X02 and X32 and X51) xor (X02 and X32 and X53) xor (X02 and X33 and X51) xor (X02 and X33 and X52) xor (X03 and X31 and X52) xor (X03 and X32 and X51) xor (X03 and X32 and X53) xor (X03 and X33 and X51) xor (X03 and X33 and X53) xor (X11 and X31 and X51) xor (X11 and X31 and X52) xor (X11 and X32 and X52) xor (X11 and X32 and X53) xor (X11 and X33 and X52) xor (X12 and X31 and X52) xor (X12 and X31 and X53) xor (X12 and X32 and X51) xor (X12 and X32 and X53) xor (X12 and X33 and X51) xor (X12 and X33 and X52) xor (X13 and X31 and X52) xor (X13 and X32 and X51) xor (X13 and X32 and X53) xor (X13 and X33 and X51) xor (X13 and X33 and X53) xor (X41 and X51) xor (X41 and X52) xor (X42 and X51) xor (X41 and X53) xor (X0_1 and X41 and X51) xor (X0_1 and X41 and X52) xor (X0_1 and X42 and X52) xor (X0_1 and X42 and X53) xor (X0_1 and X43 and X52) xor (X02 and X41 and X52) xor (X02 and X41 and X53) xor (X02 and X42 and X51) xor (X02 and X42 and X53) xor (X02 and X43 and X51) xor (X02 and X43 and X52) xor (X03 and X41 and X52) xor (X03 and X42 and X51) xor (X03 and X42 and X53) xor (X03 and X43 and X51) xor (X03 and X43 and X53) xor (X11 and X41 and X51) xor (X11 and X41 and X52) xor (X11 and X42 and X52) xor (X11 and X42 and X53) xor (X11 and X43 and X52) xor (X12 and X41 and X52) xor (X12 and X41 and X53) xor (X12 and X42 and X51) xor (X12 and X42 and X53) xor (X12 and X43 and X51) xor (X12 and X43 and X52) xor (X13 and X41 and X52) xor (X13 and X42 and X51) xor (X13 and X42 and X53) xor (X13 and X43 and X51) xor (X13 and X43 and X53) xor (X31 and X41 and X51) xor (X31 and X41 and X52) xor (X31 and X42 and X52) xor (X31 and X42 and X53) xor (X31 and X43 and X52) xor (X32 and X41 and X52) xor (X32 and X41 and X53) xor (X32 and X42 and X51) xor (X32 and X42 and X53) xor (X32 and X43 and X51) xor (X32 and X43 and X52) xor (X33 and X41 and X52) xor (X33 and X42 and X51) xor (X33 and X42 and X53) xor (X33 and X43 and X51) xor (X33 and X43 and X53) xor (X0_1 and X61) xor (X0_1 and X62) xor (X02 and X61) xor (X0_1 and X63) xor (X11 and X61) xor (X11 and X62) xor (X12 and X61) xor (X11 and X63) xor (X21 and X61) xor (X21 and X62) xor (X22 and X61) xor (X21 and X63) xor (X0_1 and X21 and X61) xor (X0_1 and X21 and X62) xor (X0_1 and X22 and X62) xor (X0_1 and X22 and X63) xor (X0_1 and X23 and X62) xor (X02 and X21 and X62) xor (X02 and X21 and X63) xor (X02 and X22 and X61) xor (X02 and X22 and X63) xor (X02 and X23 and X61) xor (X02 and X23 and X62) xor (X03 and X21 and X62) xor (X03 and X22 and X61) xor (X03 and X22 and X63) xor (X03 and X23 and X61) xor (X03 and X23 and X63) xor (X0_1 and X41 and X61) xor (X0_1 and X41 and X62) xor (X0_1 and X42 and X62) xor (X0_1 and X42 and X63) xor (X0_1 and X43 and X62) xor (X02 and X41 and X62) xor (X02 and X41 and X63) xor (X02 and X42 and X61) xor (X02 and X42 and X63) xor (X02 and X43 and X61) xor (X02 and X43 and X62) xor (X03 and X41 and X62) xor (X03 and X42 and X61) xor (X03 and X42 and X63) xor (X03 and X43 and X61) xor (X03 and X43 and X63) xor (X11 and X41 and X61) xor (X11 and X41 and X62) xor (X11 and X42 and X62) xor (X11 and X42 and X63) xor (X11 and X43 and X62) xor (X12 and X41 and X62) xor (X12 and X41 and X63) xor (X12 and X42 and X61) xor (X12 and X42 and X63) xor (X12 and X43 and X61) xor (X12 and X43 and X62) xor (X13 and X41 and X62) xor (X13 and X42 and X61) xor (X13 and X42 and X63) xor (X13 and X43 and X61) xor (X13 and X43 and X63) xor (X21 and X41 and X61) xor (X21 and X41 and X62) xor (X21 and X42 and X62) xor (X21 and X42 and X63) xor (X21 and X43 and X62) xor (X22 and X41 and X62) xor (X22 and X41 and X63) xor (X22 and X42 and X61) xor (X22 and X42 and X63) xor (X22 and X43 and X61) xor (X22 and X43 and X62) xor (X23 and X41 and X62) xor (X23 and X42 and X61) xor (X23 and X42 and X63) xor (X23 and X43 and X61) xor (X23 and X43 and X63) xor (X0_1 and X51 and X61) xor (X0_1 and X51 and X62) xor (X0_1 and X52 and X62) xor (X0_1 and X52 and X63) xor (X0_1 and X53 and X62) xor (X02 and X51 and X62) xor (X02 and X51 and X63) xor (X02 and X52 and X61) xor (X02 and X52 and X63) xor (X02 and X53 and X61) xor (X02 and X53 and X62) xor (X03 and X51 and X62) xor (X03 and X52 and X61) xor (X03 and X52 and X63) xor (X03 and X53 and X61) xor (X03 and X53 and X63) xor (X11 and X51 and X61) xor (X11 and X51 and X62) xor (X11 and X52 and X62) xor (X11 and X52 and X63) xor (X11 and X53 and X62) xor (X12 and X51 and X62) xor (X12 and X51 and X63) xor (X12 and X52 and X61) xor (X12 and X52 and X63) xor (X12 and X53 and X61) xor (X12 and X53 and X62) xor (X13 and X51 and X62) xor (X13 and X52 and X61) xor (X13 and X52 and X63) xor (X13 and X53 and X61) xor (X13 and X53 and X63) xor (X21 and X51 and X61) xor (X21 and X51 and X62) xor (X21 and X52 and X62) xor (X21 and X52 and X63) xor (X21 and X53 and X62) xor (X22 and X51 and X62) xor (X22 and X51 and X63) xor (X22 and X52 and X61) xor (X22 and X52 and X63) xor (X22 and X53 and X61) xor (X22 and X53 and X62) xor (X23 and X51 and X62) xor (X23 and X52 and X61) xor (X23 and X52 and X63) xor (X23 and X53 and X61) xor (X23 and X53 and X63) xor (X31 and X51 and X61) xor (X31 and X51 and X62) xor (X31 and X52 and X62) xor (X31 and X52 and X63) xor (X31 and X53 and X62) xor (X32 and X51 and X62) xor (X32 and X51 and X63) xor (X32 and X52 and X61) xor (X32 and X52 and X63) xor (X32 and X53 and X61) xor (X32 and X53 and X62) xor (X33 and X51 and X62) xor (X33 and X52 and X61) xor (X33 and X52 and X63) xor (X33 and X53 and X61) xor (X33 and X53 and X63) xor (X41 and X51 and X61) xor (X41 and X51 and X62) xor (X41 and X52 and X62) xor (X41 and X52 and X63) xor (X41 and X53 and X62) xor (X42 and X51 and X62) xor (X42 and X51 and X63) xor (X42 and X52 and X61) xor (X42 and X52 and X63) xor (X42 and X53 and X61) xor (X42 and X53 and X62) xor (X43 and X51 and X62) xor (X43 and X52 and X61) xor (X43 and X52 and X63) xor (X43 and X53 and X61) xor (X43 and X53 and X63) xor (X71) xor (X0_1 and X11 and X71) xor (X0_1 and X11 and X72) xor (X0_1 and X12 and X72) xor (X0_1 and X12 and X73) xor (X0_1 and X13 and X72) xor (X02 and X11 and X72) xor (X02 and X11 and X73) xor (X02 and X12 and X71) xor (X02 and X12 and X73) xor (X02 and X13 and X71) xor (X02 and X13 and X72) xor (X03 and X11 and X72) xor (X03 and X12 and X71) xor (X03 and X12 and X73) xor (X03 and X13 and X71) xor (X03 and X13 and X73) xor (X21 and X71) xor (X21 and X72) xor (X22 and X71) xor (X21 and X73) xor (X0_1 and X21 and X71) xor (X0_1 and X21 and X72) xor (X0_1 and X22 and X72) xor (X0_1 and X22 and X73) xor (X0_1 and X23 and X72) xor (X02 and X21 and X72) xor (X02 and X21 and X73) xor (X02 and X22 and X71) xor (X02 and X22 and X73) xor (X02 and X23 and X71) xor (X02 and X23 and X72) xor (X03 and X21 and X72) xor (X03 and X22 and X71) xor (X03 and X22 and X73) xor (X03 and X23 and X71) xor (X03 and X23 and X73) xor (X41 and X71) xor (X41 and X72) xor (X42 and X71) xor (X41 and X73) xor (X21 and X41 and X71) xor (X21 and X41 and X72) xor (X21 and X42 and X72) xor (X21 and X42 and X73) xor (X21 and X43 and X72) xor (X22 and X41 and X72) xor (X22 and X41 and X73) xor (X22 and X42 and X71) xor (X22 and X42 and X73) xor (X22 and X43 and X71) xor (X22 and X43 and X72) xor (X23 and X41 and X72) xor (X23 and X42 and X71) xor (X23 and X42 and X73) xor (X23 and X43 and X71) xor (X23 and X43 and X73) xor (X21 and X51 and X71) xor (X21 and X51 and X72) xor (X21 and X52 and X72) xor (X21 and X52 and X73) xor (X21 and X53 and X72) xor (X22 and X51 and X72) xor (X22 and X51 and X73) xor (X22 and X52 and X71) xor (X22 and X52 and X73) xor (X22 and X53 and X71) xor (X22 and X53 and X72) xor (X23 and X51 and X72) xor (X23 and X52 and X71) xor (X23 and X52 and X73) xor (X23 and X53 and X71) xor (X23 and X53 and X73) xor (X61 and X71) xor (X61 and X72) xor (X62 and X71) xor (X61 and X73) xor (X0_1 and X61 and X71) xor (X0_1 and X61 and X72) xor (X0_1 and X62 and X72) xor (X0_1 and X62 and X73) xor (X0_1 and X63 and X72) xor (X02 and X61 and X72) xor (X02 and X61 and X73) xor (X02 and X62 and X71) xor (X02 and X62 and X73) xor (X02 and X63 and X71) xor (X02 and X63 and X72) xor (X03 and X61 and X72) xor (X03 and X62 and X71) xor (X03 and X62 and X73) xor (X03 and X63 and X71) xor (X03 and X63 and X73) xor (X31 and X61 and X71) xor (X31 and X61 and X72) xor (X31 and X62 and X72) xor (X31 and X62 and X73) xor (X31 and X63 and X72) xor (X32 and X61 and X72) xor (X32 and X61 and X73) xor (X32 and X62 and X71) xor (X32 and X62 and X73) xor (X32 and X63 and X71) xor (X32 and X63 and X72) xor (X33 and X61 and X72) xor (X33 and X62 and X71) xor (X33 and X62 and X73) xor (X33 and X63 and X71) xor (X33 and X63 and X73) xor (X41 and X61 and X71) xor (X41 and X61 and X72) xor (X41 and X62 and X72) xor (X41 and X62 and X73) xor (X41 and X63 and X72) xor (X42 and X61 and X72) xor (X42 and X61 and X73) xor (X42 and X62 and X71) xor (X42 and X62 and X73) xor (X42 and X63 and X71) xor (X42 and X63 and X72) xor (X43 and X61 and X72) xor (X43 and X62 and X71) xor (X43 and X62 and X73) xor (X43 and X63 and X71) xor (X43 and X63 and X73) xor (X51 and X61 and X71) xor (X51 and X61 and X72) xor (X51 and X62 and X72) xor (X51 and X62 and X73) xor (X51 and X63 and X72) xor (X52 and X61 and X72) xor (X52 and X61 and X73) xor (X52 and X62 and X71) xor (X52 and X62 and X73) xor (X52 and X63 and X71) xor (X52 and X63 and X72) xor (X53 and X61 and X72) xor (X53 and X62 and X71) xor (X53 and X62 and X73) xor (X53 and X63 and X71) xor (X53 and X63 and X73));
    F72  <= ((X12) xor (X12 and X32) xor (X10 and X33) xor (X12 and X33) xor (X13 and X32) xor (X00 and X10 and X33) xor (X00 and X12 and X30) xor (X00 and X12 and X32) xor (X00 and X12 and X33) xor (X00 and X13 and X30) xor (X00 and X13 and X32) xor (X02 and X10 and X32) xor (X02 and X10 and X33) xor (X02 and X13 and X30) xor (X02 and X13 and X33) xor (X03 and X10 and X30) xor (X03 and X10 and X32) xor (X03 and X10 and X33) xor (X03 and X12 and X30) xor (X03 and X12 and X32) xor (X03 and X13 and X32) xor (X22 and X32) xor (X20 and X33) xor (X22 and X33) xor (X23 and X32) xor (X42) xor (X12 and X42) xor (X10 and X43) xor (X12 and X43) xor (X13 and X42) xor (X22 and X42) xor (X20 and X43) xor (X22 and X43) xor (X23 and X42) xor (X00 and X20 and X43) xor (X00 and X22 and X40) xor (X00 and X22 and X42) xor (X00 and X22 and X43) xor (X00 and X23 and X40) xor (X00 and X23 and X42) xor (X02 and X20 and X42) xor (X02 and X20 and X43) xor (X02 and X23 and X40) xor (X02 and X23 and X43) xor (X03 and X20 and X40) xor (X03 and X20 and X42) xor (X03 and X20 and X43) xor (X03 and X22 and X40) xor (X03 and X22 and X42) xor (X03 and X23 and X42) xor (X32 and X42) xor (X30 and X43) xor (X32 and X43) xor (X33 and X42) xor (X02 and X52) xor (X00 and X53) xor (X02 and X53) xor (X03 and X52) xor (X22 and X52) xor (X20 and X53) xor (X22 and X53) xor (X23 and X52) xor (X00 and X20 and X53) xor (X00 and X22 and X50) xor (X00 and X22 and X52) xor (X00 and X22 and X53) xor (X00 and X23 and X50) xor (X00 and X23 and X52) xor (X02 and X20 and X52) xor (X02 and X20 and X53) xor (X02 and X23 and X50) xor (X02 and X23 and X53) xor (X03 and X20 and X50) xor (X03 and X20 and X52) xor (X03 and X20 and X53) xor (X03 and X22 and X50) xor (X03 and X22 and X52) xor (X03 and X23 and X52) xor (X32 and X52) xor (X30 and X53) xor (X32 and X53) xor (X33 and X52) xor (X00 and X30 and X53) xor (X00 and X32 and X50) xor (X00 and X32 and X52) xor (X00 and X32 and X53) xor (X00 and X33 and X50) xor (X00 and X33 and X52) xor (X02 and X30 and X52) xor (X02 and X30 and X53) xor (X02 and X33 and X50) xor (X02 and X33 and X53) xor (X03 and X30 and X50) xor (X03 and X30 and X52) xor (X03 and X30 and X53) xor (X03 and X32 and X50) xor (X03 and X32 and X52) xor (X03 and X33 and X52) xor (X10 and X30 and X53) xor (X10 and X32 and X50) xor (X10 and X32 and X52) xor (X10 and X32 and X53) xor (X10 and X33 and X50) xor (X10 and X33 and X52) xor (X12 and X30 and X52) xor (X12 and X30 and X53) xor (X12 and X33 and X50) xor (X12 and X33 and X53) xor (X13 and X30 and X50) xor (X13 and X30 and X52) xor (X13 and X30 and X53) xor (X13 and X32 and X50) xor (X13 and X32 and X52) xor (X13 and X33 and X52) xor (X42 and X52) xor (X40 and X53) xor (X42 and X53) xor (X43 and X52) xor (X00 and X40 and X53) xor (X00 and X42 and X50) xor (X00 and X42 and X52) xor (X00 and X42 and X53) xor (X00 and X43 and X50) xor (X00 and X43 and X52) xor (X02 and X40 and X52) xor (X02 and X40 and X53) xor (X02 and X43 and X50) xor (X02 and X43 and X53) xor (X03 and X40 and X50) xor (X03 and X40 and X52) xor (X03 and X40 and X53) xor (X03 and X42 and X50) xor (X03 and X42 and X52) xor (X03 and X43 and X52) xor (X10 and X40 and X53) xor (X10 and X42 and X50) xor (X10 and X42 and X52) xor (X10 and X42 and X53) xor (X10 and X43 and X50) xor (X10 and X43 and X52) xor (X12 and X40 and X52) xor (X12 and X40 and X53) xor (X12 and X43 and X50) xor (X12 and X43 and X53) xor (X13 and X40 and X50) xor (X13 and X40 and X52) xor (X13 and X40 and X53) xor (X13 and X42 and X50) xor (X13 and X42 and X52) xor (X13 and X43 and X52) xor (X30 and X40 and X53) xor (X30 and X42 and X50) xor (X30 and X42 and X52) xor (X30 and X42 and X53) xor (X30 and X43 and X50) xor (X30 and X43 and X52) xor (X32 and X40 and X52) xor (X32 and X40 and X53) xor (X32 and X43 and X50) xor (X32 and X43 and X53) xor (X33 and X40 and X50) xor (X33 and X40 and X52) xor (X33 and X40 and X53) xor (X33 and X42 and X50) xor (X33 and X42 and X52) xor (X33 and X43 and X52) xor (X02 and X62) xor (X00 and X63) xor (X02 and X63) xor (X03 and X62) xor (X12 and X62) xor (X10 and X63) xor (X12 and X63) xor (X13 and X62) xor (X22 and X62) xor (X20 and X63) xor (X22 and X63) xor (X23 and X62) xor (X00 and X20 and X63) xor (X00 and X22 and X60) xor (X00 and X22 and X62) xor (X00 and X22 and X63) xor (X00 and X23 and X60) xor (X00 and X23 and X62) xor (X02 and X20 and X62) xor (X02 and X20 and X63) xor (X02 and X23 and X60) xor (X02 and X23 and X63) xor (X03 and X20 and X60) xor (X03 and X20 and X62) xor (X03 and X20 and X63) xor (X03 and X22 and X60) xor (X03 and X22 and X62) xor (X03 and X23 and X62) xor (X00 and X40 and X63) xor (X00 and X42 and X60) xor (X00 and X42 and X62) xor (X00 and X42 and X63) xor (X00 and X43 and X60) xor (X00 and X43 and X62) xor (X02 and X40 and X62) xor (X02 and X40 and X63) xor (X02 and X43 and X60) xor (X02 and X43 and X63) xor (X03 and X40 and X60) xor (X03 and X40 and X62) xor (X03 and X40 and X63) xor (X03 and X42 and X60) xor (X03 and X42 and X62) xor (X03 and X43 and X62) xor (X10 and X40 and X63) xor (X10 and X42 and X60) xor (X10 and X42 and X62) xor (X10 and X42 and X63) xor (X10 and X43 and X60) xor (X10 and X43 and X62) xor (X12 and X40 and X62) xor (X12 and X40 and X63) xor (X12 and X43 and X60) xor (X12 and X43 and X63) xor (X13 and X40 and X60) xor (X13 and X40 and X62) xor (X13 and X40 and X63) xor (X13 and X42 and X60) xor (X13 and X42 and X62) xor (X13 and X43 and X62) xor (X20 and X40 and X63) xor (X20 and X42 and X60) xor (X20 and X42 and X62) xor (X20 and X42 and X63) xor (X20 and X43 and X60) xor (X20 and X43 and X62) xor (X22 and X40 and X62) xor (X22 and X40 and X63) xor (X22 and X43 and X60) xor (X22 and X43 and X63) xor (X23 and X40 and X60) xor (X23 and X40 and X62) xor (X23 and X40 and X63) xor (X23 and X42 and X60) xor (X23 and X42 and X62) xor (X23 and X43 and X62) xor (X00 and X50 and X63) xor (X00 and X52 and X60) xor (X00 and X52 and X62) xor (X00 and X52 and X63) xor (X00 and X53 and X60) xor (X00 and X53 and X62) xor (X02 and X50 and X62) xor (X02 and X50 and X63) xor (X02 and X53 and X60) xor (X02 and X53 and X63) xor (X03 and X50 and X60) xor (X03 and X50 and X62) xor (X03 and X50 and X63) xor (X03 and X52 and X60) xor (X03 and X52 and X62) xor (X03 and X53 and X62) xor (X10 and X50 and X63) xor (X10 and X52 and X60) xor (X10 and X52 and X62) xor (X10 and X52 and X63) xor (X10 and X53 and X60) xor (X10 and X53 and X62) xor (X12 and X50 and X62) xor (X12 and X50 and X63) xor (X12 and X53 and X60) xor (X12 and X53 and X63) xor (X13 and X50 and X60) xor (X13 and X50 and X62) xor (X13 and X50 and X63) xor (X13 and X52 and X60) xor (X13 and X52 and X62) xor (X13 and X53 and X62) xor (X20 and X50 and X63) xor (X20 and X52 and X60) xor (X20 and X52 and X62) xor (X20 and X52 and X63) xor (X20 and X53 and X60) xor (X20 and X53 and X62) xor (X22 and X50 and X62) xor (X22 and X50 and X63) xor (X22 and X53 and X60) xor (X22 and X53 and X63) xor (X23 and X50 and X60) xor (X23 and X50 and X62) xor (X23 and X50 and X63) xor (X23 and X52 and X60) xor (X23 and X52 and X62) xor (X23 and X53 and X62) xor (X30 and X50 and X63) xor (X30 and X52 and X60) xor (X30 and X52 and X62) xor (X30 and X52 and X63) xor (X30 and X53 and X60) xor (X30 and X53 and X62) xor (X32 and X50 and X62) xor (X32 and X50 and X63) xor (X32 and X53 and X60) xor (X32 and X53 and X63) xor (X33 and X50 and X60) xor (X33 and X50 and X62) xor (X33 and X50 and X63) xor (X33 and X52 and X60) xor (X33 and X52 and X62) xor (X33 and X53 and X62) xor (X40 and X50 and X63) xor (X40 and X52 and X60) xor (X40 and X52 and X62) xor (X40 and X52 and X63) xor (X40 and X53 and X60) xor (X40 and X53 and X62) xor (X42 and X50 and X62) xor (X42 and X50 and X63) xor (X42 and X53 and X60) xor (X42 and X53 and X63) xor (X43 and X50 and X60) xor (X43 and X50 and X62) xor (X43 and X50 and X63) xor (X43 and X52 and X60) xor (X43 and X52 and X62) xor (X43 and X53 and X62) xor (X72) xor (X00 and X10 and X73) xor (X00 and X12 and X70) xor (X00 and X12 and X72) xor (X00 and X12 and X73) xor (X00 and X13 and X70) xor (X00 and X13 and X72) xor (X02 and X10 and X72) xor (X02 and X10 and X73) xor (X02 and X13 and X70) xor (X02 and X13 and X73) xor (X03 and X10 and X70) xor (X03 and X10 and X72) xor (X03 and X10 and X73) xor (X03 and X12 and X70) xor (X03 and X12 and X72) xor (X03 and X13 and X72) xor (X22 and X72) xor (X20 and X73) xor (X22 and X73) xor (X23 and X72) xor (X00 and X20 and X73) xor (X00 and X22 and X70) xor (X00 and X22 and X72) xor (X00 and X22 and X73) xor (X00 and X23 and X70) xor (X00 and X23 and X72) xor (X02 and X20 and X72) xor (X02 and X20 and X73) xor (X02 and X23 and X70) xor (X02 and X23 and X73) xor (X03 and X20 and X70) xor (X03 and X20 and X72) xor (X03 and X20 and X73) xor (X03 and X22 and X70) xor (X03 and X22 and X72) xor (X03 and X23 and X72) xor (X42 and X72) xor (X40 and X73) xor (X42 and X73) xor (X43 and X72) xor (X20 and X40 and X73) xor (X20 and X42 and X70) xor (X20 and X42 and X72) xor (X20 and X42 and X73) xor (X20 and X43 and X70) xor (X20 and X43 and X72) xor (X22 and X40 and X72) xor (X22 and X40 and X73) xor (X22 and X43 and X70) xor (X22 and X43 and X73) xor (X23 and X40 and X70) xor (X23 and X40 and X72) xor (X23 and X40 and X73) xor (X23 and X42 and X70) xor (X23 and X42 and X72) xor (X23 and X43 and X72) xor (X20 and X50 and X73) xor (X20 and X52 and X70) xor (X20 and X52 and X72) xor (X20 and X52 and X73) xor (X20 and X53 and X70) xor (X20 and X53 and X72) xor (X22 and X50 and X72) xor (X22 and X50 and X73) xor (X22 and X53 and X70) xor (X22 and X53 and X73) xor (X23 and X50 and X70) xor (X23 and X50 and X72) xor (X23 and X50 and X73) xor (X23 and X52 and X70) xor (X23 and X52 and X72) xor (X23 and X53 and X72) xor (X62 and X72) xor (X60 and X73) xor (X62 and X73) xor (X63 and X72) xor (X00 and X60 and X73) xor (X00 and X62 and X70) xor (X00 and X62 and X72) xor (X00 and X62 and X73) xor (X00 and X63 and X70) xor (X00 and X63 and X72) xor (X02 and X60 and X72) xor (X02 and X60 and X73) xor (X02 and X63 and X70) xor (X02 and X63 and X73) xor (X03 and X60 and X70) xor (X03 and X60 and X72) xor (X03 and X60 and X73) xor (X03 and X62 and X70) xor (X03 and X62 and X72) xor (X03 and X63 and X72) xor (X30 and X60 and X73) xor (X30 and X62 and X70) xor (X30 and X62 and X72) xor (X30 and X62 and X73) xor (X30 and X63 and X70) xor (X30 and X63 and X72) xor (X32 and X60 and X72) xor (X32 and X60 and X73) xor (X32 and X63 and X70) xor (X32 and X63 and X73) xor (X33 and X60 and X70) xor (X33 and X60 and X72) xor (X33 and X60 and X73) xor (X33 and X62 and X70) xor (X33 and X62 and X72) xor (X33 and X63 and X72) xor (X40 and X60 and X73) xor (X40 and X62 and X70) xor (X40 and X62 and X72) xor (X40 and X62 and X73) xor (X40 and X63 and X70) xor (X40 and X63 and X72) xor (X42 and X60 and X72) xor (X42 and X60 and X73) xor (X42 and X63 and X70) xor (X42 and X63 and X73) xor (X43 and X60 and X70) xor (X43 and X60 and X72) xor (X43 and X60 and X73) xor (X43 and X62 and X70) xor (X43 and X62 and X72) xor (X43 and X63 and X72) xor (X50 and X60 and X73) xor (X50 and X62 and X70) xor (X50 and X62 and X72) xor (X50 and X62 and X73) xor (X50 and X63 and X70) xor (X50 and X63 and X72) xor (X52 and X60 and X72) xor (X52 and X60 and X73) xor (X52 and X63 and X70) xor (X52 and X63 and X73) xor (X53 and X60 and X70) xor (X53 and X60 and X72) xor (X53 and X60 and X73) xor (X53 and X62 and X70) xor (X53 and X62 and X72) xor (X53 and X63 and X72));
    F73  <= ((X13) xor (X13 and X33) xor (X13 and X30) xor (X13 and X31) xor (X11 and X30) xor (X00 and X10 and X31) xor (X00 and X11 and X30) xor (X00 and X11 and X33) xor (X00 and X13 and X31) xor (X00 and X13 and X33) xor (X0_1 and X10 and X31) xor (X0_1 and X10 and X33) xor (X0_1 and X11 and X33) xor (X0_1 and X13 and X30) xor (X0_1 and X13 and X31) xor (X0_1 and X13 and X33) xor (X03 and X10 and X31) xor (X03 and X11 and X30) xor (X03 and X11 and X31) xor (X03 and X11 and X33) xor (X03 and X13 and X30) xor (X23 and X33) xor (X23 and X30) xor (X23 and X31) xor (X21 and X30) xor (X43) xor (X13 and X43) xor (X13 and X40) xor (X13 and X41) xor (X11 and X40) xor (X23 and X43) xor (X23 and X40) xor (X23 and X41) xor (X21 and X40) xor (X00 and X20 and X41) xor (X00 and X21 and X40) xor (X00 and X21 and X43) xor (X00 and X23 and X41) xor (X00 and X23 and X43) xor (X0_1 and X20 and X41) xor (X0_1 and X20 and X43) xor (X0_1 and X21 and X43) xor (X0_1 and X23 and X40) xor (X0_1 and X23 and X41) xor (X0_1 and X23 and X43) xor (X03 and X20 and X41) xor (X03 and X21 and X40) xor (X03 and X21 and X41) xor (X03 and X21 and X43) xor (X03 and X23 and X40) xor (X33 and X43) xor (X33 and X40) xor (X33 and X41) xor (X31 and X40) xor (X03 and X53) xor (X03 and X50) xor (X03 and X51) xor (X0_1 and X50) xor (X23 and X53) xor (X23 and X50) xor (X23 and X51) xor (X21 and X50) xor (X00 and X20 and X51) xor (X00 and X21 and X50) xor (X00 and X21 and X53) xor (X00 and X23 and X51) xor (X00 and X23 and X53) xor (X0_1 and X20 and X51) xor (X0_1 and X20 and X53) xor (X0_1 and X21 and X53) xor (X0_1 and X23 and X50) xor (X0_1 and X23 and X51) xor (X0_1 and X23 and X53) xor (X03 and X20 and X51) xor (X03 and X21 and X50) xor (X03 and X21 and X51) xor (X03 and X21 and X53) xor (X03 and X23 and X50) xor (X33 and X53) xor (X33 and X50) xor (X33 and X51) xor (X31 and X50) xor (X00 and X30 and X51) xor (X00 and X31 and X50) xor (X00 and X31 and X53) xor (X00 and X33 and X51) xor (X00 and X33 and X53) xor (X0_1 and X30 and X51) xor (X0_1 and X30 and X53) xor (X0_1 and X31 and X53) xor (X0_1 and X33 and X50) xor (X0_1 and X33 and X51) xor (X0_1 and X33 and X53) xor (X03 and X30 and X51) xor (X03 and X31 and X50) xor (X03 and X31 and X51) xor (X03 and X31 and X53) xor (X03 and X33 and X50) xor (X10 and X30 and X51) xor (X10 and X31 and X50) xor (X10 and X31 and X53) xor (X10 and X33 and X51) xor (X10 and X33 and X53) xor (X11 and X30 and X51) xor (X11 and X30 and X53) xor (X11 and X31 and X53) xor (X11 and X33 and X50) xor (X11 and X33 and X51) xor (X11 and X33 and X53) xor (X13 and X30 and X51) xor (X13 and X31 and X50) xor (X13 and X31 and X51) xor (X13 and X31 and X53) xor (X13 and X33 and X50) xor (X43 and X53) xor (X43 and X50) xor (X43 and X51) xor (X41 and X50) xor (X00 and X40 and X51) xor (X00 and X41 and X50) xor (X00 and X41 and X53) xor (X00 and X43 and X51) xor (X00 and X43 and X53) xor (X0_1 and X40 and X51) xor (X0_1 and X40 and X53) xor (X0_1 and X41 and X53) xor (X0_1 and X43 and X50) xor (X0_1 and X43 and X51) xor (X0_1 and X43 and X53) xor (X03 and X40 and X51) xor (X03 and X41 and X50) xor (X03 and X41 and X51) xor (X03 and X41 and X53) xor (X03 and X43 and X50) xor (X10 and X40 and X51) xor (X10 and X41 and X50) xor (X10 and X41 and X53) xor (X10 and X43 and X51) xor (X10 and X43 and X53) xor (X11 and X40 and X51) xor (X11 and X40 and X53) xor (X11 and X41 and X53) xor (X11 and X43 and X50) xor (X11 and X43 and X51) xor (X11 and X43 and X53) xor (X13 and X40 and X51) xor (X13 and X41 and X50) xor (X13 and X41 and X51) xor (X13 and X41 and X53) xor (X13 and X43 and X50) xor (X30 and X40 and X51) xor (X30 and X41 and X50) xor (X30 and X41 and X53) xor (X30 and X43 and X51) xor (X30 and X43 and X53) xor (X31 and X40 and X51) xor (X31 and X40 and X53) xor (X31 and X41 and X53) xor (X31 and X43 and X50) xor (X31 and X43 and X51) xor (X31 and X43 and X53) xor (X33 and X40 and X51) xor (X33 and X41 and X50) xor (X33 and X41 and X51) xor (X33 and X41 and X53) xor (X33 and X43 and X50) xor (X03 and X63) xor (X03 and X60) xor (X03 and X61) xor (X0_1 and X60) xor (X13 and X63) xor (X13 and X60) xor (X13 and X61) xor (X11 and X60) xor (X23 and X63) xor (X23 and X60) xor (X23 and X61) xor (X21 and X60) xor (X00 and X20 and X61) xor (X00 and X21 and X60) xor (X00 and X21 and X63) xor (X00 and X23 and X61) xor (X00 and X23 and X63) xor (X0_1 and X20 and X61) xor (X0_1 and X20 and X63) xor (X0_1 and X21 and X63) xor (X0_1 and X23 and X60) xor (X0_1 and X23 and X61) xor (X0_1 and X23 and X63) xor (X03 and X20 and X61) xor (X03 and X21 and X60) xor (X03 and X21 and X61) xor (X03 and X21 and X63) xor (X03 and X23 and X60) xor (X00 and X40 and X61) xor (X00 and X41 and X60) xor (X00 and X41 and X63) xor (X00 and X43 and X61) xor (X00 and X43 and X63) xor (X0_1 and X40 and X61) xor (X0_1 and X40 and X63) xor (X0_1 and X41 and X63) xor (X0_1 and X43 and X60) xor (X0_1 and X43 and X61) xor (X0_1 and X43 and X63) xor (X03 and X40 and X61) xor (X03 and X41 and X60) xor (X03 and X41 and X61) xor (X03 and X41 and X63) xor (X03 and X43 and X60) xor (X10 and X40 and X61) xor (X10 and X41 and X60) xor (X10 and X41 and X63) xor (X10 and X43 and X61) xor (X10 and X43 and X63) xor (X11 and X40 and X61) xor (X11 and X40 and X63) xor (X11 and X41 and X63) xor (X11 and X43 and X60) xor (X11 and X43 and X61) xor (X11 and X43 and X63) xor (X13 and X40 and X61) xor (X13 and X41 and X60) xor (X13 and X41 and X61) xor (X13 and X41 and X63) xor (X13 and X43 and X60) xor (X20 and X40 and X61) xor (X20 and X41 and X60) xor (X20 and X41 and X63) xor (X20 and X43 and X61) xor (X20 and X43 and X63) xor (X21 and X40 and X61) xor (X21 and X40 and X63) xor (X21 and X41 and X63) xor (X21 and X43 and X60) xor (X21 and X43 and X61) xor (X21 and X43 and X63) xor (X23 and X40 and X61) xor (X23 and X41 and X60) xor (X23 and X41 and X61) xor (X23 and X41 and X63) xor (X23 and X43 and X60) xor (X00 and X50 and X61) xor (X00 and X51 and X60) xor (X00 and X51 and X63) xor (X00 and X53 and X61) xor (X00 and X53 and X63) xor (X0_1 and X50 and X61) xor (X0_1 and X50 and X63) xor (X0_1 and X51 and X63) xor (X0_1 and X53 and X60) xor (X0_1 and X53 and X61) xor (X0_1 and X53 and X63) xor (X03 and X50 and X61) xor (X03 and X51 and X60) xor (X03 and X51 and X61) xor (X03 and X51 and X63) xor (X03 and X53 and X60) xor (X10 and X50 and X61) xor (X10 and X51 and X60) xor (X10 and X51 and X63) xor (X10 and X53 and X61) xor (X10 and X53 and X63) xor (X11 and X50 and X61) xor (X11 and X50 and X63) xor (X11 and X51 and X63) xor (X11 and X53 and X60) xor (X11 and X53 and X61) xor (X11 and X53 and X63) xor (X13 and X50 and X61) xor (X13 and X51 and X60) xor (X13 and X51 and X61) xor (X13 and X51 and X63) xor (X13 and X53 and X60) xor (X20 and X50 and X61) xor (X20 and X51 and X60) xor (X20 and X51 and X63) xor (X20 and X53 and X61) xor (X20 and X53 and X63) xor (X21 and X50 and X61) xor (X21 and X50 and X63) xor (X21 and X51 and X63) xor (X21 and X53 and X60) xor (X21 and X53 and X61) xor (X21 and X53 and X63) xor (X23 and X50 and X61) xor (X23 and X51 and X60) xor (X23 and X51 and X61) xor (X23 and X51 and X63) xor (X23 and X53 and X60) xor (X30 and X50 and X61) xor (X30 and X51 and X60) xor (X30 and X51 and X63) xor (X30 and X53 and X61) xor (X30 and X53 and X63) xor (X31 and X50 and X61) xor (X31 and X50 and X63) xor (X31 and X51 and X63) xor (X31 and X53 and X60) xor (X31 and X53 and X61) xor (X31 and X53 and X63) xor (X33 and X50 and X61) xor (X33 and X51 and X60) xor (X33 and X51 and X61) xor (X33 and X51 and X63) xor (X33 and X53 and X60) xor (X40 and X50 and X61) xor (X40 and X51 and X60) xor (X40 and X51 and X63) xor (X40 and X53 and X61) xor (X40 and X53 and X63) xor (X41 and X50 and X61) xor (X41 and X50 and X63) xor (X41 and X51 and X63) xor (X41 and X53 and X60) xor (X41 and X53 and X61) xor (X41 and X53 and X63) xor (X43 and X50 and X61) xor (X43 and X51 and X60) xor (X43 and X51 and X61) xor (X43 and X51 and X63) xor (X43 and X53 and X60) xor (X73) xor (X00 and X10 and X71) xor (X00 and X11 and X70) xor (X00 and X11 and X73) xor (X00 and X13 and X71) xor (X00 and X13 and X73) xor (X0_1 and X10 and X71) xor (X0_1 and X10 and X73) xor (X0_1 and X11 and X73) xor (X0_1 and X13 and X70) xor (X0_1 and X13 and X71) xor (X0_1 and X13 and X73) xor (X03 and X10 and X71) xor (X03 and X11 and X70) xor (X03 and X11 and X71) xor (X03 and X11 and X73) xor (X03 and X13 and X70) xor (X23 and X73) xor (X23 and X70) xor (X23 and X71) xor (X21 and X70) xor (X00 and X20 and X71) xor (X00 and X21 and X70) xor (X00 and X21 and X73) xor (X00 and X23 and X71) xor (X00 and X23 and X73) xor (X0_1 and X20 and X71) xor (X0_1 and X20 and X73) xor (X0_1 and X21 and X73) xor (X0_1 and X23 and X70) xor (X0_1 and X23 and X71) xor (X0_1 and X23 and X73) xor (X03 and X20 and X71) xor (X03 and X21 and X70) xor (X03 and X21 and X71) xor (X03 and X21 and X73) xor (X03 and X23 and X70) xor (X43 and X73) xor (X43 and X70) xor (X43 and X71) xor (X41 and X70) xor (X20 and X40 and X71) xor (X20 and X41 and X70) xor (X20 and X41 and X73) xor (X20 and X43 and X71) xor (X20 and X43 and X73) xor (X21 and X40 and X71) xor (X21 and X40 and X73) xor (X21 and X41 and X73) xor (X21 and X43 and X70) xor (X21 and X43 and X71) xor (X21 and X43 and X73) xor (X23 and X40 and X71) xor (X23 and X41 and X70) xor (X23 and X41 and X71) xor (X23 and X41 and X73) xor (X23 and X43 and X70) xor (X20 and X50 and X71) xor (X20 and X51 and X70) xor (X20 and X51 and X73) xor (X20 and X53 and X71) xor (X20 and X53 and X73) xor (X21 and X50 and X71) xor (X21 and X50 and X73) xor (X21 and X51 and X73) xor (X21 and X53 and X70) xor (X21 and X53 and X71) xor (X21 and X53 and X73) xor (X23 and X50 and X71) xor (X23 and X51 and X70) xor (X23 and X51 and X71) xor (X23 and X51 and X73) xor (X23 and X53 and X70) xor (X63 and X73) xor (X63 and X70) xor (X63 and X71) xor (X61 and X70) xor (X00 and X60 and X71) xor (X00 and X61 and X70) xor (X00 and X61 and X73) xor (X00 and X63 and X71) xor (X00 and X63 and X73) xor (X0_1 and X60 and X71) xor (X0_1 and X60 and X73) xor (X0_1 and X61 and X73) xor (X0_1 and X63 and X70) xor (X0_1 and X63 and X71) xor (X0_1 and X63 and X73) xor (X03 and X60 and X71) xor (X03 and X61 and X70) xor (X03 and X61 and X71) xor (X03 and X61 and X73) xor (X03 and X63 and X70) xor (X30 and X60 and X71) xor (X30 and X61 and X70) xor (X30 and X61 and X73) xor (X30 and X63 and X71) xor (X30 and X63 and X73) xor (X31 and X60 and X71) xor (X31 and X60 and X73) xor (X31 and X61 and X73) xor (X31 and X63 and X70) xor (X31 and X63 and X71) xor (X31 and X63 and X73) xor (X33 and X60 and X71) xor (X33 and X61 and X70) xor (X33 and X61 and X71) xor (X33 and X61 and X73) xor (X33 and X63 and X70) xor (X40 and X60 and X71) xor (X40 and X61 and X70) xor (X40 and X61 and X73) xor (X40 and X63 and X71) xor (X40 and X63 and X73) xor (X41 and X60 and X71) xor (X41 and X60 and X73) xor (X41 and X61 and X73) xor (X41 and X63 and X70) xor (X41 and X63 and X71) xor (X41 and X63 and X73) xor (X43 and X60 and X71) xor (X43 and X61 and X70) xor (X43 and X61 and X71) xor (X43 and X61 and X73) xor (X43 and X63 and X70) xor (X50 and X60 and X71) xor (X50 and X61 and X70) xor (X50 and X61 and X73) xor (X50 and X63 and X71) xor (X50 and X63 and X73) xor (X51 and X60 and X71) xor (X51 and X60 and X73) xor (X51 and X61 and X73) xor (X51 and X63 and X70) xor (X51 and X63 and X71) xor (X51 and X63 and X73) xor (X53 and X60 and X71) xor (X53 and X61 and X70) xor (X53 and X61 and X71) xor (X53 and X61 and X73) xor (X53 and X63 and X70));
end Behavioral;
